magic
tech sky130A
magscale 1 2
timestamp 1733308831
<< viali >>
rect 1593 7497 1627 7531
rect 4169 7497 4203 7531
rect 5825 7497 5859 7531
rect 7941 7497 7975 7531
rect 10057 7497 10091 7531
rect 12173 7497 12207 7531
rect 14289 7497 14323 7531
rect 16865 7497 16899 7531
rect 18889 7497 18923 7531
rect 21005 7497 21039 7531
rect 23581 7497 23615 7531
rect 24869 7497 24903 7531
rect 27169 7497 27203 7531
rect 27537 7497 27571 7531
rect 29101 7497 29135 7531
rect 31217 7497 31251 7531
rect 33333 7497 33367 7531
rect 35449 7497 35483 7531
rect 37565 7497 37599 7531
rect 37933 7497 37967 7531
rect 40049 7497 40083 7531
rect 41797 7497 41831 7531
rect 43453 7497 43487 7531
rect 3893 7429 3927 7463
rect 18429 7429 18463 7463
rect 20545 7429 20579 7463
rect 20913 7429 20947 7463
rect 27077 7429 27111 7463
rect 33241 7429 33275 7463
rect 1501 7361 1535 7395
rect 5733 7361 5767 7395
rect 7849 7361 7883 7395
rect 9965 7361 9999 7395
rect 12081 7361 12115 7395
rect 14197 7361 14231 7395
rect 16773 7361 16807 7395
rect 19073 7361 19107 7395
rect 21189 7361 21223 7395
rect 22845 7361 22879 7395
rect 23305 7361 23339 7395
rect 23489 7361 23523 7395
rect 24777 7361 24811 7395
rect 27721 7361 27755 7395
rect 29009 7361 29043 7395
rect 31125 7361 31159 7395
rect 35357 7361 35391 7395
rect 37473 7361 37507 7395
rect 38117 7361 38151 7395
rect 39957 7361 39991 7395
rect 41705 7361 41739 7395
rect 43177 7361 43211 7395
rect 23121 7225 23155 7259
rect 18521 7157 18555 7191
rect 23029 6749 23063 6783
rect 22845 6613 22879 6647
rect 16589 5865 16623 5899
rect 24869 5865 24903 5899
rect 16129 5661 16163 5695
rect 16405 5661 16439 5695
rect 25053 5661 25087 5695
rect 25513 3689 25547 3723
rect 27813 3689 27847 3723
rect 29193 3689 29227 3723
rect 33609 3689 33643 3723
rect 17417 3621 17451 3655
rect 23029 3621 23063 3655
rect 24685 3621 24719 3655
rect 26617 3621 26651 3655
rect 28365 3621 28399 3655
rect 17049 3485 17083 3519
rect 17601 3485 17635 3519
rect 18705 3485 18739 3519
rect 18981 3485 19015 3519
rect 19533 3485 19567 3519
rect 19901 3485 19935 3519
rect 20177 3485 20211 3519
rect 20821 3485 20855 3519
rect 21097 3485 21131 3519
rect 21373 3485 21407 3519
rect 21649 3485 21683 3519
rect 21925 3485 21959 3519
rect 22201 3485 22235 3519
rect 22661 3485 22695 3519
rect 23213 3485 23247 3519
rect 23489 3485 23523 3519
rect 24593 3485 24627 3519
rect 24869 3485 24903 3519
rect 25421 3485 25455 3519
rect 25697 3485 25731 3519
rect 25973 3485 26007 3519
rect 26249 3485 26283 3519
rect 26525 3485 26559 3519
rect 26801 3485 26835 3519
rect 27077 3485 27111 3519
rect 27445 3485 27479 3519
rect 27997 3485 28031 3519
rect 28273 3485 28307 3519
rect 28549 3485 28583 3519
rect 28825 3485 28859 3519
rect 29377 3485 29411 3519
rect 32965 3417 32999 3451
rect 33517 3417 33551 3451
rect 16865 3349 16899 3383
rect 18521 3349 18555 3383
rect 18797 3349 18831 3383
rect 19349 3349 19383 3383
rect 19717 3349 19751 3383
rect 19993 3349 20027 3383
rect 20637 3349 20671 3383
rect 20913 3349 20947 3383
rect 21189 3349 21223 3383
rect 21465 3349 21499 3383
rect 21741 3349 21775 3383
rect 22017 3349 22051 3383
rect 22477 3349 22511 3383
rect 23305 3349 23339 3383
rect 24409 3349 24443 3383
rect 25237 3349 25271 3383
rect 25789 3349 25823 3383
rect 26065 3349 26099 3383
rect 26341 3349 26375 3383
rect 26893 3349 26927 3383
rect 27261 3349 27295 3383
rect 28089 3349 28123 3383
rect 28641 3349 28675 3383
rect 33057 3349 33091 3383
rect 9321 3145 9355 3179
rect 13921 3145 13955 3179
rect 14565 3145 14599 3179
rect 14841 3145 14875 3179
rect 19165 3145 19199 3179
rect 24041 3145 24075 3179
rect 31585 3145 31619 3179
rect 33977 3145 34011 3179
rect 35081 3145 35115 3179
rect 35449 3145 35483 3179
rect 38117 3145 38151 3179
rect 20729 3077 20763 3111
rect 21281 3077 21315 3111
rect 22201 3077 22235 3111
rect 22753 3077 22787 3111
rect 23305 3077 23339 3111
rect 24685 3077 24719 3111
rect 27629 3077 27663 3111
rect 29285 3077 29319 3111
rect 29837 3077 29871 3111
rect 30941 3077 30975 3111
rect 34437 3077 34471 3111
rect 34989 3077 35023 3111
rect 9137 3009 9171 3043
rect 13737 3009 13771 3043
rect 14381 3009 14415 3043
rect 14657 3009 14691 3043
rect 14933 3009 14967 3043
rect 15393 3009 15427 3043
rect 15669 3009 15703 3043
rect 15945 3009 15979 3043
rect 16221 3009 16255 3043
rect 16497 3009 16531 3043
rect 16957 3009 16991 3043
rect 17049 3009 17083 3043
rect 17509 3009 17543 3043
rect 17785 3009 17819 3043
rect 17877 3009 17911 3043
rect 18153 3009 18187 3043
rect 18613 3009 18647 3043
rect 18705 3009 18739 3043
rect 18981 3009 19015 3043
rect 19257 3009 19291 3043
rect 19625 3009 19659 3043
rect 20177 3009 20211 3043
rect 22017 3009 22051 3043
rect 23949 3009 23983 3043
rect 24225 3009 24259 3043
rect 24501 3009 24535 3043
rect 25237 3009 25271 3043
rect 25789 3009 25823 3043
rect 26341 3009 26375 3043
rect 27077 3009 27111 3043
rect 28181 3009 28215 3043
rect 28733 3009 28767 3043
rect 30389 3009 30423 3043
rect 31493 3009 31527 3043
rect 32781 3009 32815 3043
rect 33333 3009 33367 3043
rect 33885 3009 33919 3043
rect 35357 3009 35391 3043
rect 35817 3009 35851 3043
rect 36093 3009 36127 3043
rect 36185 3009 36219 3043
rect 38025 3009 38059 3043
rect 38301 3009 38335 3043
rect 39129 3009 39163 3043
rect 39405 3009 39439 3043
rect 16773 2873 16807 2907
rect 17601 2873 17635 2907
rect 18337 2873 18371 2907
rect 18429 2873 18463 2907
rect 19441 2873 19475 2907
rect 19809 2873 19843 2907
rect 35633 2873 35667 2907
rect 37841 2873 37875 2907
rect 15117 2805 15151 2839
rect 15209 2805 15243 2839
rect 15485 2805 15519 2839
rect 15761 2805 15795 2839
rect 16037 2805 16071 2839
rect 16313 2805 16347 2839
rect 17233 2805 17267 2839
rect 17325 2805 17359 2839
rect 18061 2805 18095 2839
rect 18889 2805 18923 2839
rect 20269 2805 20303 2839
rect 20821 2805 20855 2839
rect 21373 2805 21407 2839
rect 21833 2805 21867 2839
rect 22293 2805 22327 2839
rect 22845 2805 22879 2839
rect 23397 2805 23431 2839
rect 23765 2805 23799 2839
rect 24317 2805 24351 2839
rect 24777 2805 24811 2839
rect 25329 2805 25363 2839
rect 25881 2805 25915 2839
rect 26433 2805 26467 2839
rect 27169 2805 27203 2839
rect 27721 2805 27755 2839
rect 28273 2805 28307 2839
rect 28825 2805 28859 2839
rect 29377 2805 29411 2839
rect 29929 2805 29963 2839
rect 30481 2805 30515 2839
rect 31033 2805 31067 2839
rect 32321 2805 32355 2839
rect 32873 2805 32907 2839
rect 33425 2805 33459 2839
rect 34529 2805 34563 2839
rect 35909 2805 35943 2839
rect 36369 2805 36403 2839
rect 38945 2805 38979 2839
rect 39221 2805 39255 2839
rect 5641 2601 5675 2635
rect 8769 2601 8803 2635
rect 9413 2601 9447 2635
rect 9965 2601 9999 2635
rect 10241 2601 10275 2635
rect 11069 2601 11103 2635
rect 13921 2601 13955 2635
rect 14105 2601 14139 2635
rect 17233 2601 17267 2635
rect 25697 2601 25731 2635
rect 26617 2601 26651 2635
rect 27721 2601 27755 2635
rect 28825 2601 28859 2635
rect 29193 2601 29227 2635
rect 30849 2601 30883 2635
rect 31769 2601 31803 2635
rect 32873 2601 32907 2635
rect 34345 2601 34379 2635
rect 36737 2601 36771 2635
rect 36829 2601 36863 2635
rect 39221 2601 39255 2635
rect 40141 2601 40175 2635
rect 40417 2601 40451 2635
rect 41245 2601 41279 2635
rect 42809 2601 42843 2635
rect 4813 2533 4847 2567
rect 6193 2533 6227 2567
rect 7113 2533 7147 2567
rect 9137 2533 9171 2567
rect 9505 2533 9539 2567
rect 11713 2533 11747 2567
rect 11989 2533 12023 2567
rect 12265 2533 12299 2567
rect 12541 2533 12575 2567
rect 13093 2533 13127 2567
rect 13461 2533 13495 2567
rect 17141 2533 17175 2567
rect 18061 2533 18095 2567
rect 19257 2533 19291 2567
rect 21833 2533 21867 2567
rect 28365 2533 28399 2567
rect 30389 2533 30423 2567
rect 35541 2533 35575 2567
rect 36093 2533 36127 2567
rect 37289 2533 37323 2567
rect 39129 2533 39163 2567
rect 39865 2533 39899 2567
rect 40693 2533 40727 2567
rect 40969 2533 41003 2567
rect 33609 2465 33643 2499
rect 4629 2397 4663 2431
rect 4905 2397 4939 2431
rect 5181 2397 5215 2431
rect 5457 2397 5491 2431
rect 5733 2397 5767 2431
rect 6009 2397 6043 2431
rect 6377 2397 6411 2431
rect 6653 2397 6687 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 8033 2397 8067 2431
rect 8309 2397 8343 2431
rect 8585 2397 8619 2431
rect 8953 2397 8987 2431
rect 9229 2397 9263 2431
rect 9689 2397 9723 2431
rect 9781 2397 9815 2431
rect 10057 2397 10091 2431
rect 10333 2397 10367 2431
rect 10609 2397 10643 2431
rect 10885 2397 10919 2431
rect 11161 2397 11195 2431
rect 11529 2397 11563 2431
rect 11805 2397 11839 2431
rect 12081 2397 12115 2431
rect 12357 2397 12391 2431
rect 12633 2397 12667 2431
rect 12909 2397 12943 2431
rect 13185 2397 13219 2431
rect 13645 2397 13679 2431
rect 13737 2397 13771 2431
rect 14289 2397 14323 2431
rect 14933 2397 14967 2431
rect 15209 2397 15243 2431
rect 15485 2397 15519 2431
rect 15761 2397 15795 2431
rect 16037 2397 16071 2431
rect 16313 2397 16347 2431
rect 16681 2397 16715 2431
rect 16957 2397 16991 2431
rect 17417 2397 17451 2431
rect 17693 2397 17727 2431
rect 17785 2397 17819 2431
rect 18245 2397 18279 2431
rect 18521 2397 18555 2431
rect 19441 2397 19475 2431
rect 19625 2397 19659 2431
rect 20177 2397 20211 2431
rect 20729 2397 20763 2431
rect 21281 2397 21315 2431
rect 22017 2397 22051 2431
rect 22201 2397 22235 2431
rect 22753 2397 22787 2431
rect 23305 2397 23339 2431
rect 23857 2397 23891 2431
rect 24501 2397 24535 2431
rect 25053 2397 25087 2431
rect 26157 2397 26191 2431
rect 26801 2397 26835 2431
rect 27077 2397 27111 2431
rect 28181 2397 28215 2431
rect 28733 2397 28767 2431
rect 29377 2397 29411 2431
rect 29653 2397 29687 2431
rect 30205 2397 30239 2431
rect 31309 2397 31343 2431
rect 31953 2397 31987 2431
rect 34529 2397 34563 2431
rect 35909 2397 35943 2431
rect 36277 2397 36311 2431
rect 36553 2397 36587 2431
rect 37013 2397 37047 2431
rect 37473 2397 37507 2431
rect 37565 2397 37599 2431
rect 37841 2397 37875 2431
rect 38117 2397 38151 2431
rect 38393 2397 38427 2431
rect 38669 2397 38703 2431
rect 38945 2397 38979 2431
rect 39405 2397 39439 2431
rect 39681 2397 39715 2431
rect 40049 2397 40083 2431
rect 40325 2397 40359 2431
rect 40601 2397 40635 2431
rect 40877 2397 40911 2431
rect 41153 2397 41187 2431
rect 41429 2397 41463 2431
rect 42993 2397 43027 2431
rect 18705 2329 18739 2363
rect 19073 2329 19107 2363
rect 19993 2329 20027 2363
rect 20545 2329 20579 2363
rect 21097 2329 21131 2363
rect 21649 2329 21683 2363
rect 25605 2329 25639 2363
rect 27629 2329 27663 2363
rect 30757 2329 30791 2363
rect 32229 2329 32263 2363
rect 32781 2329 32815 2363
rect 33333 2329 33367 2363
rect 33885 2329 33919 2363
rect 34805 2329 34839 2363
rect 35357 2329 35391 2363
rect 5089 2261 5123 2295
rect 5365 2261 5399 2295
rect 5917 2261 5951 2295
rect 6561 2261 6595 2295
rect 6837 2261 6871 2295
rect 7389 2261 7423 2295
rect 7665 2261 7699 2295
rect 7941 2261 7975 2295
rect 8217 2261 8251 2295
rect 8493 2261 8527 2295
rect 10517 2261 10551 2295
rect 10793 2261 10827 2295
rect 11345 2261 11379 2295
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 14657 2261 14691 2295
rect 15117 2261 15151 2295
rect 15393 2261 15427 2295
rect 15669 2261 15703 2295
rect 15945 2261 15979 2295
rect 16221 2261 16255 2295
rect 16497 2261 16531 2295
rect 16865 2261 16899 2295
rect 17509 2261 17543 2295
rect 17969 2261 18003 2295
rect 18337 2261 18371 2295
rect 22293 2261 22327 2295
rect 22845 2261 22879 2295
rect 23581 2261 23615 2295
rect 23949 2261 23983 2295
rect 24593 2261 24627 2295
rect 25145 2261 25179 2295
rect 26249 2261 26283 2295
rect 27169 2261 27203 2295
rect 29745 2261 29779 2295
rect 31401 2261 31435 2295
rect 32321 2261 32355 2295
rect 33977 2261 34011 2295
rect 34897 2261 34931 2295
rect 36369 2261 36403 2295
rect 37749 2261 37783 2295
rect 38025 2261 38059 2295
rect 38301 2261 38335 2295
rect 38577 2261 38611 2295
rect 38853 2261 38887 2295
rect 39497 2261 39531 2295
<< metal1 >>
rect 22186 7760 22192 7812
rect 22244 7800 22250 7812
rect 31386 7800 31392 7812
rect 22244 7772 31392 7800
rect 22244 7760 22250 7772
rect 31386 7760 31392 7772
rect 31444 7760 31450 7812
rect 19058 7692 19064 7744
rect 19116 7732 19122 7744
rect 35894 7732 35900 7744
rect 19116 7704 35900 7732
rect 19116 7692 19122 7704
rect 35894 7692 35900 7704
rect 35952 7692 35958 7744
rect 1104 7642 44040 7664
rect 1104 7590 11644 7642
rect 11696 7590 11708 7642
rect 11760 7590 11772 7642
rect 11824 7590 11836 7642
rect 11888 7590 11900 7642
rect 11952 7590 22338 7642
rect 22390 7590 22402 7642
rect 22454 7590 22466 7642
rect 22518 7590 22530 7642
rect 22582 7590 22594 7642
rect 22646 7590 33032 7642
rect 33084 7590 33096 7642
rect 33148 7590 33160 7642
rect 33212 7590 33224 7642
rect 33276 7590 33288 7642
rect 33340 7590 43726 7642
rect 43778 7590 43790 7642
rect 43842 7590 43854 7642
rect 43906 7590 43918 7642
rect 43970 7590 43982 7642
rect 44034 7590 44040 7642
rect 1104 7568 44040 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 1360 7500 1593 7528
rect 1360 7488 1366 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 4157 7531 4215 7537
rect 4157 7528 4169 7531
rect 3844 7500 4169 7528
rect 3844 7488 3850 7500
rect 4157 7497 4169 7500
rect 4203 7497 4215 7531
rect 4157 7491 4215 7497
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5592 7500 5825 7528
rect 5592 7488 5598 7500
rect 5813 7497 5825 7500
rect 5859 7497 5871 7531
rect 5813 7491 5871 7497
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 7708 7500 7941 7528
rect 7708 7488 7714 7500
rect 7929 7497 7941 7500
rect 7975 7497 7987 7531
rect 7929 7491 7987 7497
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 10045 7531 10103 7537
rect 10045 7528 10057 7531
rect 9824 7500 10057 7528
rect 9824 7488 9830 7500
rect 10045 7497 10057 7500
rect 10091 7497 10103 7531
rect 10045 7491 10103 7497
rect 12158 7488 12164 7540
rect 12216 7488 12222 7540
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14277 7531 14335 7537
rect 14277 7528 14289 7531
rect 14056 7500 14289 7528
rect 14056 7488 14062 7500
rect 14277 7497 14289 7500
rect 14323 7497 14335 7531
rect 14277 7491 14335 7497
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 16632 7500 16865 7528
rect 16632 7488 16638 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 16853 7491 16911 7497
rect 18877 7531 18935 7537
rect 18877 7497 18889 7531
rect 18923 7497 18935 7531
rect 20993 7531 21051 7537
rect 20993 7528 21005 7531
rect 18877 7491 18935 7497
rect 20548 7500 21005 7528
rect 3881 7463 3939 7469
rect 3881 7429 3893 7463
rect 3927 7460 3939 7463
rect 18417 7463 18475 7469
rect 3927 7432 17264 7460
rect 3927 7429 3939 7432
rect 3881 7423 3939 7429
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 4062 7392 4068 7404
rect 1535 7364 4068 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 5718 7352 5724 7404
rect 5776 7352 5782 7404
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 7852 7188 7880 7355
rect 9968 7256 9996 7355
rect 12084 7324 12112 7355
rect 14182 7352 14188 7404
rect 14240 7352 14246 7404
rect 16758 7352 16764 7404
rect 16816 7352 16822 7404
rect 17236 7392 17264 7432
rect 18417 7429 18429 7463
rect 18463 7460 18475 7463
rect 18892 7460 18920 7491
rect 20548 7469 20576 7500
rect 20993 7497 21005 7500
rect 21039 7497 21051 7531
rect 20993 7491 21051 7497
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 21140 7500 22094 7528
rect 21140 7488 21146 7500
rect 18463 7432 18920 7460
rect 20533 7463 20591 7469
rect 18463 7429 18475 7432
rect 18417 7423 18475 7429
rect 20533 7429 20545 7463
rect 20579 7429 20591 7463
rect 20533 7423 20591 7429
rect 20714 7420 20720 7472
rect 20772 7460 20778 7472
rect 20901 7463 20959 7469
rect 20901 7460 20913 7463
rect 20772 7432 20913 7460
rect 20772 7420 20778 7432
rect 20901 7429 20913 7432
rect 20947 7429 20959 7463
rect 22066 7460 22094 7500
rect 22830 7488 22836 7540
rect 22888 7528 22894 7540
rect 23569 7531 23627 7537
rect 23569 7528 23581 7531
rect 22888 7500 23581 7528
rect 22888 7488 22894 7500
rect 23569 7497 23581 7500
rect 23615 7497 23627 7531
rect 23569 7491 23627 7497
rect 24670 7488 24676 7540
rect 24728 7528 24734 7540
rect 24857 7531 24915 7537
rect 24857 7528 24869 7531
rect 24728 7500 24869 7528
rect 24728 7488 24734 7500
rect 24857 7497 24869 7500
rect 24903 7497 24915 7531
rect 24857 7491 24915 7497
rect 26694 7488 26700 7540
rect 26752 7528 26758 7540
rect 27157 7531 27215 7537
rect 27157 7528 27169 7531
rect 26752 7500 27169 7528
rect 26752 7488 26758 7500
rect 27157 7497 27169 7500
rect 27203 7497 27215 7531
rect 27157 7491 27215 7497
rect 27525 7531 27583 7537
rect 27525 7497 27537 7531
rect 27571 7497 27583 7531
rect 27525 7491 27583 7497
rect 27065 7463 27123 7469
rect 22066 7432 26924 7460
rect 20901 7423 20959 7429
rect 26896 7404 26924 7432
rect 27065 7429 27077 7463
rect 27111 7460 27123 7463
rect 27540 7460 27568 7491
rect 28902 7488 28908 7540
rect 28960 7528 28966 7540
rect 29089 7531 29147 7537
rect 29089 7528 29101 7531
rect 28960 7500 29101 7528
rect 28960 7488 28966 7500
rect 29089 7497 29101 7500
rect 29135 7497 29147 7531
rect 29089 7491 29147 7497
rect 30926 7488 30932 7540
rect 30984 7528 30990 7540
rect 31205 7531 31263 7537
rect 31205 7528 31217 7531
rect 30984 7500 31217 7528
rect 30984 7488 30990 7500
rect 31205 7497 31217 7500
rect 31251 7497 31263 7531
rect 31205 7491 31263 7497
rect 32950 7488 32956 7540
rect 33008 7528 33014 7540
rect 33321 7531 33379 7537
rect 33321 7528 33333 7531
rect 33008 7500 33333 7528
rect 33008 7488 33014 7500
rect 33321 7497 33333 7500
rect 33367 7497 33379 7531
rect 33321 7491 33379 7497
rect 35158 7488 35164 7540
rect 35216 7528 35222 7540
rect 35437 7531 35495 7537
rect 35437 7528 35449 7531
rect 35216 7500 35449 7528
rect 35216 7488 35222 7500
rect 35437 7497 35449 7500
rect 35483 7497 35495 7531
rect 35437 7491 35495 7497
rect 37274 7488 37280 7540
rect 37332 7528 37338 7540
rect 37553 7531 37611 7537
rect 37553 7528 37565 7531
rect 37332 7500 37565 7528
rect 37332 7488 37338 7500
rect 37553 7497 37565 7500
rect 37599 7497 37611 7531
rect 37553 7491 37611 7497
rect 37921 7531 37979 7537
rect 37921 7497 37933 7531
rect 37967 7497 37979 7531
rect 37921 7491 37979 7497
rect 33229 7463 33287 7469
rect 27111 7432 27568 7460
rect 27614 7432 31892 7460
rect 27111 7429 27123 7432
rect 27065 7423 27123 7429
rect 18598 7392 18604 7404
rect 17236 7364 18604 7392
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 19058 7352 19064 7404
rect 19116 7352 19122 7404
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7392 21235 7395
rect 21910 7392 21916 7404
rect 21223 7364 21916 7392
rect 21223 7361 21235 7364
rect 21177 7355 21235 7361
rect 21910 7352 21916 7364
rect 21968 7352 21974 7404
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7392 22891 7395
rect 23293 7395 23351 7401
rect 23293 7392 23305 7395
rect 22879 7364 23305 7392
rect 22879 7361 22891 7364
rect 22833 7355 22891 7361
rect 23293 7361 23305 7364
rect 23339 7392 23351 7395
rect 23382 7392 23388 7404
rect 23339 7364 23388 7392
rect 23339 7361 23351 7364
rect 23293 7355 23351 7361
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 23474 7352 23480 7404
rect 23532 7352 23538 7404
rect 24765 7395 24823 7401
rect 24765 7361 24777 7395
rect 24811 7392 24823 7395
rect 24854 7392 24860 7404
rect 24811 7364 24860 7392
rect 24811 7361 24823 7364
rect 24765 7355 24823 7361
rect 24854 7352 24860 7364
rect 24912 7352 24918 7404
rect 26878 7352 26884 7404
rect 26936 7352 26942 7404
rect 27614 7324 27642 7432
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 12084 7296 27642 7324
rect 27724 7324 27752 7355
rect 28994 7352 29000 7404
rect 29052 7352 29058 7404
rect 31113 7395 31171 7401
rect 31113 7361 31125 7395
rect 31159 7392 31171 7395
rect 31754 7392 31760 7404
rect 31159 7364 31760 7392
rect 31159 7361 31171 7364
rect 31113 7355 31171 7361
rect 31754 7352 31760 7364
rect 31812 7352 31818 7404
rect 31864 7392 31892 7432
rect 33229 7429 33241 7463
rect 33275 7460 33287 7463
rect 37936 7460 37964 7491
rect 39666 7488 39672 7540
rect 39724 7528 39730 7540
rect 40037 7531 40095 7537
rect 40037 7528 40049 7531
rect 39724 7500 40049 7528
rect 39724 7488 39730 7500
rect 40037 7497 40049 7500
rect 40083 7497 40095 7531
rect 40037 7491 40095 7497
rect 41506 7488 41512 7540
rect 41564 7528 41570 7540
rect 41785 7531 41843 7537
rect 41785 7528 41797 7531
rect 41564 7500 41797 7528
rect 41564 7488 41570 7500
rect 41785 7497 41797 7500
rect 41831 7497 41843 7531
rect 41785 7491 41843 7497
rect 43441 7531 43499 7537
rect 43441 7497 43453 7531
rect 43487 7528 43499 7531
rect 43622 7528 43628 7540
rect 43487 7500 43628 7528
rect 43487 7497 43499 7500
rect 43441 7491 43499 7497
rect 43622 7488 43628 7500
rect 43680 7488 43686 7540
rect 33275 7432 37964 7460
rect 33275 7429 33287 7432
rect 33229 7423 33287 7429
rect 31864 7364 34468 7392
rect 34330 7324 34336 7336
rect 27724 7296 34336 7324
rect 34330 7284 34336 7296
rect 34388 7284 34394 7336
rect 34440 7324 34468 7364
rect 35342 7352 35348 7404
rect 35400 7352 35406 7404
rect 37461 7395 37519 7401
rect 37461 7361 37473 7395
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 38105 7395 38163 7401
rect 38105 7361 38117 7395
rect 38151 7361 38163 7395
rect 38105 7355 38163 7361
rect 39945 7395 40003 7401
rect 39945 7361 39957 7395
rect 39991 7392 40003 7395
rect 40218 7392 40224 7404
rect 39991 7364 40224 7392
rect 39991 7361 40003 7364
rect 39945 7355 40003 7361
rect 35526 7324 35532 7336
rect 34440 7296 35532 7324
rect 35526 7284 35532 7296
rect 35584 7284 35590 7336
rect 22186 7256 22192 7268
rect 9968 7228 22192 7256
rect 22186 7216 22192 7228
rect 22244 7216 22250 7268
rect 23109 7259 23167 7265
rect 23109 7256 23121 7259
rect 22664 7228 23121 7256
rect 17310 7188 17316 7200
rect 7852 7160 17316 7188
rect 17310 7148 17316 7160
rect 17368 7148 17374 7200
rect 18230 7148 18236 7200
rect 18288 7188 18294 7200
rect 18509 7191 18567 7197
rect 18509 7188 18521 7191
rect 18288 7160 18521 7188
rect 18288 7148 18294 7160
rect 18509 7157 18521 7160
rect 18555 7157 18567 7191
rect 18509 7151 18567 7157
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 22664 7188 22692 7228
rect 23109 7225 23121 7228
rect 23155 7225 23167 7259
rect 37476 7256 37504 7355
rect 38120 7324 38148 7355
rect 40218 7352 40224 7364
rect 40276 7352 40282 7404
rect 41690 7352 41696 7404
rect 41748 7352 41754 7404
rect 43162 7352 43168 7404
rect 43220 7352 43226 7404
rect 40494 7324 40500 7336
rect 38120 7296 40500 7324
rect 40494 7284 40500 7296
rect 40552 7284 40558 7336
rect 40034 7256 40040 7268
rect 37476 7228 40040 7256
rect 23109 7219 23167 7225
rect 40034 7216 40040 7228
rect 40092 7216 40098 7268
rect 18656 7160 22692 7188
rect 18656 7148 18662 7160
rect 1104 7098 43884 7120
rect 1104 7046 6297 7098
rect 6349 7046 6361 7098
rect 6413 7046 6425 7098
rect 6477 7046 6489 7098
rect 6541 7046 6553 7098
rect 6605 7046 16991 7098
rect 17043 7046 17055 7098
rect 17107 7046 17119 7098
rect 17171 7046 17183 7098
rect 17235 7046 17247 7098
rect 17299 7046 27685 7098
rect 27737 7046 27749 7098
rect 27801 7046 27813 7098
rect 27865 7046 27877 7098
rect 27929 7046 27941 7098
rect 27993 7046 38379 7098
rect 38431 7046 38443 7098
rect 38495 7046 38507 7098
rect 38559 7046 38571 7098
rect 38623 7046 38635 7098
rect 38687 7046 43884 7098
rect 1104 7024 43884 7046
rect 17310 6944 17316 6996
rect 17368 6984 17374 6996
rect 21082 6984 21088 6996
rect 17368 6956 21088 6984
rect 17368 6944 17374 6956
rect 21082 6944 21088 6956
rect 21140 6944 21146 6996
rect 23382 6944 23388 6996
rect 23440 6984 23446 6996
rect 36722 6984 36728 6996
rect 23440 6956 36728 6984
rect 23440 6944 23446 6956
rect 36722 6944 36728 6956
rect 36780 6944 36786 6996
rect 26878 6876 26884 6928
rect 26936 6916 26942 6928
rect 34422 6916 34428 6928
rect 26936 6888 34428 6916
rect 26936 6876 26942 6888
rect 34422 6876 34428 6888
rect 34480 6876 34486 6928
rect 23014 6740 23020 6792
rect 23072 6740 23078 6792
rect 23474 6740 23480 6792
rect 23532 6740 23538 6792
rect 22833 6647 22891 6653
rect 22833 6613 22845 6647
rect 22879 6644 22891 6647
rect 23492 6644 23520 6740
rect 22879 6616 23520 6644
rect 22879 6613 22891 6616
rect 22833 6607 22891 6613
rect 1104 6554 44040 6576
rect 1104 6502 11644 6554
rect 11696 6502 11708 6554
rect 11760 6502 11772 6554
rect 11824 6502 11836 6554
rect 11888 6502 11900 6554
rect 11952 6502 22338 6554
rect 22390 6502 22402 6554
rect 22454 6502 22466 6554
rect 22518 6502 22530 6554
rect 22582 6502 22594 6554
rect 22646 6502 33032 6554
rect 33084 6502 33096 6554
rect 33148 6502 33160 6554
rect 33212 6502 33224 6554
rect 33276 6502 33288 6554
rect 33340 6502 43726 6554
rect 43778 6502 43790 6554
rect 43842 6502 43854 6554
rect 43906 6502 43918 6554
rect 43970 6502 43982 6554
rect 44034 6502 44040 6554
rect 1104 6480 44040 6502
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 35802 6236 35808 6248
rect 5776 6208 35808 6236
rect 5776 6196 5782 6208
rect 35802 6196 35808 6208
rect 35860 6196 35866 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 33594 6168 33600 6180
rect 4120 6140 33600 6168
rect 4120 6128 4126 6140
rect 33594 6128 33600 6140
rect 33652 6128 33658 6180
rect 1104 6010 43884 6032
rect 1104 5958 6297 6010
rect 6349 5958 6361 6010
rect 6413 5958 6425 6010
rect 6477 5958 6489 6010
rect 6541 5958 6553 6010
rect 6605 5958 16991 6010
rect 17043 5958 17055 6010
rect 17107 5958 17119 6010
rect 17171 5958 17183 6010
rect 17235 5958 17247 6010
rect 17299 5958 27685 6010
rect 27737 5958 27749 6010
rect 27801 5958 27813 6010
rect 27865 5958 27877 6010
rect 27929 5958 27941 6010
rect 27993 5958 38379 6010
rect 38431 5958 38443 6010
rect 38495 5958 38507 6010
rect 38559 5958 38571 6010
rect 38623 5958 38635 6010
rect 38687 5958 43884 6010
rect 1104 5936 43884 5958
rect 16577 5899 16635 5905
rect 16577 5865 16589 5899
rect 16623 5896 16635 5899
rect 16758 5896 16764 5908
rect 16623 5868 16764 5896
rect 16623 5865 16635 5868
rect 16577 5859 16635 5865
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 24854 5856 24860 5908
rect 24912 5856 24918 5908
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5692 16175 5695
rect 16393 5695 16451 5701
rect 16393 5692 16405 5695
rect 16163 5664 16405 5692
rect 16163 5661 16175 5664
rect 16117 5655 16175 5661
rect 16393 5661 16405 5664
rect 16439 5692 16451 5695
rect 16482 5692 16488 5704
rect 16439 5664 16488 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 25041 5695 25099 5701
rect 25041 5661 25053 5695
rect 25087 5692 25099 5695
rect 38930 5692 38936 5704
rect 25087 5664 38936 5692
rect 25087 5661 25099 5664
rect 25041 5655 25099 5661
rect 38930 5652 38936 5664
rect 38988 5652 38994 5704
rect 35894 5516 35900 5568
rect 35952 5556 35958 5568
rect 38010 5556 38016 5568
rect 35952 5528 38016 5556
rect 35952 5516 35958 5528
rect 38010 5516 38016 5528
rect 38068 5516 38074 5568
rect 1104 5466 44040 5488
rect 1104 5414 11644 5466
rect 11696 5414 11708 5466
rect 11760 5414 11772 5466
rect 11824 5414 11836 5466
rect 11888 5414 11900 5466
rect 11952 5414 22338 5466
rect 22390 5414 22402 5466
rect 22454 5414 22466 5466
rect 22518 5414 22530 5466
rect 22582 5414 22594 5466
rect 22646 5414 33032 5466
rect 33084 5414 33096 5466
rect 33148 5414 33160 5466
rect 33212 5414 33224 5466
rect 33276 5414 33288 5466
rect 33340 5414 43726 5466
rect 43778 5414 43790 5466
rect 43842 5414 43854 5466
rect 43906 5414 43918 5466
rect 43970 5414 43982 5466
rect 44034 5414 44040 5466
rect 1104 5392 44040 5414
rect 1104 4922 43884 4944
rect 1104 4870 6297 4922
rect 6349 4870 6361 4922
rect 6413 4870 6425 4922
rect 6477 4870 6489 4922
rect 6541 4870 6553 4922
rect 6605 4870 16991 4922
rect 17043 4870 17055 4922
rect 17107 4870 17119 4922
rect 17171 4870 17183 4922
rect 17235 4870 17247 4922
rect 17299 4870 27685 4922
rect 27737 4870 27749 4922
rect 27801 4870 27813 4922
rect 27865 4870 27877 4922
rect 27929 4870 27941 4922
rect 27993 4870 38379 4922
rect 38431 4870 38443 4922
rect 38495 4870 38507 4922
rect 38559 4870 38571 4922
rect 38623 4870 38635 4922
rect 38687 4870 43884 4922
rect 1104 4848 43884 4870
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 19426 4740 19432 4752
rect 9732 4712 19432 4740
rect 9732 4700 9738 4712
rect 19426 4700 19432 4712
rect 19484 4700 19490 4752
rect 10226 4632 10232 4684
rect 10284 4672 10290 4684
rect 28810 4672 28816 4684
rect 10284 4644 28816 4672
rect 10284 4632 10290 4644
rect 28810 4632 28816 4644
rect 28868 4632 28874 4684
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 24210 4604 24216 4616
rect 6236 4576 24216 4604
rect 6236 4564 6242 4576
rect 24210 4564 24216 4576
rect 24268 4564 24274 4616
rect 14090 4496 14096 4548
rect 14148 4536 14154 4548
rect 25958 4536 25964 4548
rect 14148 4508 25964 4536
rect 14148 4496 14154 4508
rect 25958 4496 25964 4508
rect 26016 4496 26022 4548
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 24486 4468 24492 4480
rect 8720 4440 24492 4468
rect 8720 4428 8726 4440
rect 24486 4428 24492 4440
rect 24544 4428 24550 4480
rect 1104 4378 44040 4400
rect 1104 4326 11644 4378
rect 11696 4326 11708 4378
rect 11760 4326 11772 4378
rect 11824 4326 11836 4378
rect 11888 4326 11900 4378
rect 11952 4326 22338 4378
rect 22390 4326 22402 4378
rect 22454 4326 22466 4378
rect 22518 4326 22530 4378
rect 22582 4326 22594 4378
rect 22646 4326 33032 4378
rect 33084 4326 33096 4378
rect 33148 4326 33160 4378
rect 33212 4326 33224 4378
rect 33276 4326 33288 4378
rect 33340 4326 43726 4378
rect 43778 4326 43790 4378
rect 43842 4326 43854 4378
rect 43906 4326 43918 4378
rect 43970 4326 43982 4378
rect 44034 4326 44040 4378
rect 1104 4304 44040 4326
rect 14458 4224 14464 4276
rect 14516 4264 14522 4276
rect 25498 4264 25504 4276
rect 14516 4236 25504 4264
rect 14516 4224 14522 4236
rect 25498 4224 25504 4236
rect 25556 4224 25562 4276
rect 13906 4156 13912 4208
rect 13964 4196 13970 4208
rect 33410 4196 33416 4208
rect 13964 4168 33416 4196
rect 13964 4156 13970 4168
rect 33410 4156 33416 4168
rect 33468 4156 33474 4208
rect 13906 4020 13912 4072
rect 13964 4060 13970 4072
rect 13964 4032 22094 4060
rect 13964 4020 13970 4032
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 10376 3964 21772 3992
rect 10376 3952 10382 3964
rect 21744 3936 21772 3964
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 20162 3924 20168 3936
rect 10008 3896 20168 3924
rect 10008 3884 10014 3896
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 21726 3884 21732 3936
rect 21784 3884 21790 3936
rect 22066 3924 22094 4032
rect 25406 3924 25412 3936
rect 22066 3896 25412 3924
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 26234 3884 26240 3936
rect 26292 3924 26298 3936
rect 30006 3924 30012 3936
rect 26292 3896 30012 3924
rect 26292 3884 26298 3896
rect 30006 3884 30012 3896
rect 30064 3884 30070 3936
rect 1104 3834 43884 3856
rect 1104 3782 6297 3834
rect 6349 3782 6361 3834
rect 6413 3782 6425 3834
rect 6477 3782 6489 3834
rect 6541 3782 6553 3834
rect 6605 3782 16991 3834
rect 17043 3782 17055 3834
rect 17107 3782 17119 3834
rect 17171 3782 17183 3834
rect 17235 3782 17247 3834
rect 17299 3782 27685 3834
rect 27737 3782 27749 3834
rect 27801 3782 27813 3834
rect 27865 3782 27877 3834
rect 27929 3782 27941 3834
rect 27993 3782 38379 3834
rect 38431 3782 38443 3834
rect 38495 3782 38507 3834
rect 38559 3782 38571 3834
rect 38623 3782 38635 3834
rect 38687 3782 43884 3834
rect 1104 3760 43884 3782
rect 15102 3680 15108 3732
rect 15160 3720 15166 3732
rect 25501 3723 25559 3729
rect 15160 3692 24624 3720
rect 15160 3680 15166 3692
rect 16666 3612 16672 3664
rect 16724 3652 16730 3664
rect 17405 3655 17463 3661
rect 17405 3652 17417 3655
rect 16724 3624 17417 3652
rect 16724 3612 16730 3624
rect 17405 3621 17417 3624
rect 17451 3621 17463 3655
rect 17405 3615 17463 3621
rect 23017 3655 23075 3661
rect 23017 3621 23029 3655
rect 23063 3652 23075 3655
rect 23474 3652 23480 3664
rect 23063 3624 23480 3652
rect 23063 3621 23075 3624
rect 23017 3615 23075 3621
rect 23474 3612 23480 3624
rect 23532 3612 23538 3664
rect 9306 3544 9312 3596
rect 9364 3584 9370 3596
rect 9364 3556 21680 3584
rect 9364 3544 9370 3556
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 16816 3488 17049 3516
rect 16816 3476 16822 3488
rect 17037 3485 17049 3488
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 18472 3488 18705 3516
rect 18472 3476 18478 3488
rect 18693 3485 18705 3488
rect 18739 3485 18751 3519
rect 18693 3479 18751 3485
rect 18969 3519 19027 3525
rect 18969 3485 18981 3519
rect 19015 3485 19027 3519
rect 18969 3479 19027 3485
rect 18598 3408 18604 3460
rect 18656 3448 18662 3460
rect 18984 3448 19012 3479
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19300 3488 19533 3516
rect 19300 3476 19306 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 19886 3476 19892 3528
rect 19944 3476 19950 3528
rect 20162 3476 20168 3528
rect 20220 3476 20226 3528
rect 20806 3476 20812 3528
rect 20864 3476 20870 3528
rect 21085 3519 21143 3525
rect 21085 3485 21097 3519
rect 21131 3485 21143 3519
rect 21085 3479 21143 3485
rect 18656 3420 19012 3448
rect 18656 3408 18662 3420
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 21100 3448 21128 3479
rect 21358 3476 21364 3528
rect 21416 3476 21422 3528
rect 21652 3525 21680 3556
rect 22094 3544 22100 3596
rect 22152 3584 22158 3596
rect 22152 3556 22692 3584
rect 22152 3544 22158 3556
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3485 21695 3519
rect 21637 3479 21695 3485
rect 21726 3476 21732 3528
rect 21784 3516 21790 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21784 3488 21925 3516
rect 21784 3476 21790 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 22002 3476 22008 3528
rect 22060 3516 22066 3528
rect 22664 3525 22692 3556
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 22060 3488 22201 3516
rect 22060 3476 22066 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 22649 3519 22707 3525
rect 22649 3485 22661 3519
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 23198 3476 23204 3528
rect 23256 3476 23262 3528
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3516 23535 3519
rect 23842 3516 23848 3528
rect 23523 3488 23848 3516
rect 23523 3485 23535 3488
rect 23477 3479 23535 3485
rect 23842 3476 23848 3488
rect 23900 3476 23906 3528
rect 24596 3525 24624 3692
rect 25501 3689 25513 3723
rect 25547 3720 25559 3723
rect 27062 3720 27068 3732
rect 25547 3692 27068 3720
rect 25547 3689 25559 3692
rect 25501 3683 25559 3689
rect 27062 3680 27068 3692
rect 27120 3680 27126 3732
rect 27801 3723 27859 3729
rect 27801 3689 27813 3723
rect 27847 3720 27859 3723
rect 27847 3692 28304 3720
rect 27847 3689 27859 3692
rect 27801 3683 27859 3689
rect 24673 3655 24731 3661
rect 24673 3621 24685 3655
rect 24719 3652 24731 3655
rect 25682 3652 25688 3664
rect 24719 3624 25688 3652
rect 24719 3621 24731 3624
rect 24673 3615 24731 3621
rect 25682 3612 25688 3624
rect 25740 3612 25746 3664
rect 26605 3655 26663 3661
rect 26605 3621 26617 3655
rect 26651 3652 26663 3655
rect 27982 3652 27988 3664
rect 26651 3624 27988 3652
rect 26651 3621 26663 3624
rect 26605 3615 26663 3621
rect 27982 3612 27988 3624
rect 28040 3612 28046 3664
rect 24946 3544 24952 3596
rect 25004 3584 25010 3596
rect 28276 3584 28304 3692
rect 28994 3680 29000 3732
rect 29052 3720 29058 3732
rect 29181 3723 29239 3729
rect 29181 3720 29193 3723
rect 29052 3692 29193 3720
rect 29052 3680 29058 3692
rect 29181 3689 29193 3692
rect 29227 3689 29239 3723
rect 29181 3683 29239 3689
rect 33594 3680 33600 3732
rect 33652 3680 33658 3732
rect 28353 3655 28411 3661
rect 28353 3621 28365 3655
rect 28399 3652 28411 3655
rect 29822 3652 29828 3664
rect 28399 3624 29828 3652
rect 28399 3621 28411 3624
rect 28353 3615 28411 3621
rect 29822 3612 29828 3624
rect 29880 3612 29886 3664
rect 29546 3584 29552 3596
rect 25004 3556 27108 3584
rect 28276 3556 29552 3584
rect 25004 3544 25010 3556
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 19484 3420 21128 3448
rect 21744 3420 22232 3448
rect 19484 3408 19490 3420
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 16853 3383 16911 3389
rect 16853 3380 16865 3383
rect 16356 3352 16865 3380
rect 16356 3340 16362 3352
rect 16853 3349 16865 3352
rect 16899 3349 16911 3383
rect 16853 3343 16911 3349
rect 17770 3340 17776 3392
rect 17828 3380 17834 3392
rect 18509 3383 18567 3389
rect 18509 3380 18521 3383
rect 17828 3352 18521 3380
rect 17828 3340 17834 3352
rect 18509 3349 18521 3352
rect 18555 3349 18567 3383
rect 18509 3343 18567 3349
rect 18782 3340 18788 3392
rect 18840 3340 18846 3392
rect 19334 3340 19340 3392
rect 19392 3340 19398 3392
rect 19702 3340 19708 3392
rect 19760 3340 19766 3392
rect 19978 3340 19984 3392
rect 20036 3340 20042 3392
rect 20625 3383 20683 3389
rect 20625 3349 20637 3383
rect 20671 3380 20683 3383
rect 20806 3380 20812 3392
rect 20671 3352 20812 3380
rect 20671 3349 20683 3352
rect 20625 3343 20683 3349
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 20898 3340 20904 3392
rect 20956 3340 20962 3392
rect 21174 3340 21180 3392
rect 21232 3340 21238 3392
rect 21450 3340 21456 3392
rect 21508 3340 21514 3392
rect 21744 3389 21772 3420
rect 22204 3392 22232 3420
rect 23658 3408 23664 3460
rect 23716 3448 23722 3460
rect 24872 3448 24900 3479
rect 25406 3476 25412 3528
rect 25464 3476 25470 3528
rect 25498 3476 25504 3528
rect 25556 3516 25562 3528
rect 25685 3519 25743 3525
rect 25685 3516 25697 3519
rect 25556 3488 25697 3516
rect 25556 3476 25562 3488
rect 25685 3485 25697 3488
rect 25731 3485 25743 3519
rect 25685 3479 25743 3485
rect 25958 3476 25964 3528
rect 26016 3476 26022 3528
rect 26234 3476 26240 3528
rect 26292 3476 26298 3528
rect 26510 3476 26516 3528
rect 26568 3476 26574 3528
rect 26786 3476 26792 3528
rect 26844 3476 26850 3528
rect 27080 3525 27108 3556
rect 29546 3544 29552 3556
rect 29604 3544 29610 3596
rect 27065 3519 27123 3525
rect 27065 3485 27077 3519
rect 27111 3485 27123 3519
rect 27065 3479 27123 3485
rect 27154 3476 27160 3528
rect 27212 3516 27218 3528
rect 27433 3519 27491 3525
rect 27433 3516 27445 3519
rect 27212 3488 27445 3516
rect 27212 3476 27218 3488
rect 27433 3485 27445 3488
rect 27479 3485 27491 3519
rect 27433 3479 27491 3485
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 27985 3519 28043 3525
rect 27985 3516 27997 3519
rect 27672 3488 27997 3516
rect 27672 3476 27678 3488
rect 27985 3485 27997 3488
rect 28031 3485 28043 3519
rect 27985 3479 28043 3485
rect 28258 3476 28264 3528
rect 28316 3476 28322 3528
rect 28534 3476 28540 3528
rect 28592 3476 28598 3528
rect 28810 3476 28816 3528
rect 28868 3476 28874 3528
rect 29365 3519 29423 3525
rect 29365 3485 29377 3519
rect 29411 3516 29423 3519
rect 36814 3516 36820 3528
rect 29411 3488 36820 3516
rect 29411 3485 29423 3488
rect 29365 3479 29423 3485
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 26694 3448 26700 3460
rect 23716 3420 24900 3448
rect 25792 3420 26700 3448
rect 23716 3408 23722 3420
rect 21729 3383 21787 3389
rect 21729 3349 21741 3383
rect 21775 3349 21787 3383
rect 21729 3343 21787 3349
rect 22002 3340 22008 3392
rect 22060 3340 22066 3392
rect 22186 3340 22192 3392
rect 22244 3340 22250 3392
rect 22465 3383 22523 3389
rect 22465 3349 22477 3383
rect 22511 3380 22523 3383
rect 22922 3380 22928 3392
rect 22511 3352 22928 3380
rect 22511 3349 22523 3352
rect 22465 3343 22523 3349
rect 22922 3340 22928 3352
rect 22980 3340 22986 3392
rect 23293 3383 23351 3389
rect 23293 3349 23305 3383
rect 23339 3380 23351 3383
rect 23934 3380 23940 3392
rect 23339 3352 23940 3380
rect 23339 3349 23351 3352
rect 23293 3343 23351 3349
rect 23934 3340 23940 3352
rect 23992 3340 23998 3392
rect 24394 3340 24400 3392
rect 24452 3340 24458 3392
rect 25222 3340 25228 3392
rect 25280 3340 25286 3392
rect 25792 3389 25820 3420
rect 26694 3408 26700 3420
rect 26752 3408 26758 3460
rect 28718 3448 28724 3460
rect 27264 3420 28724 3448
rect 25777 3383 25835 3389
rect 25777 3349 25789 3383
rect 25823 3349 25835 3383
rect 25777 3343 25835 3349
rect 26053 3383 26111 3389
rect 26053 3349 26065 3383
rect 26099 3380 26111 3383
rect 26142 3380 26148 3392
rect 26099 3352 26148 3380
rect 26099 3349 26111 3352
rect 26053 3343 26111 3349
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 26326 3340 26332 3392
rect 26384 3340 26390 3392
rect 26878 3340 26884 3392
rect 26936 3340 26942 3392
rect 27264 3389 27292 3420
rect 28718 3408 28724 3420
rect 28776 3408 28782 3460
rect 32030 3408 32036 3460
rect 32088 3448 32094 3460
rect 32953 3451 33011 3457
rect 32953 3448 32965 3451
rect 32088 3420 32965 3448
rect 32088 3408 32094 3420
rect 32953 3417 32965 3420
rect 32999 3417 33011 3451
rect 32953 3411 33011 3417
rect 33502 3408 33508 3460
rect 33560 3408 33566 3460
rect 27249 3383 27307 3389
rect 27249 3349 27261 3383
rect 27295 3349 27307 3383
rect 27249 3343 27307 3349
rect 28074 3340 28080 3392
rect 28132 3340 28138 3392
rect 28626 3340 28632 3392
rect 28684 3340 28690 3392
rect 32766 3340 32772 3392
rect 32824 3380 32830 3392
rect 33045 3383 33103 3389
rect 33045 3380 33057 3383
rect 32824 3352 33057 3380
rect 32824 3340 32830 3352
rect 33045 3349 33057 3352
rect 33091 3349 33103 3383
rect 33045 3343 33103 3349
rect 34974 3340 34980 3392
rect 35032 3380 35038 3392
rect 36906 3380 36912 3392
rect 35032 3352 36912 3380
rect 35032 3340 35038 3352
rect 36906 3340 36912 3352
rect 36964 3340 36970 3392
rect 1104 3290 44040 3312
rect 1104 3238 11644 3290
rect 11696 3238 11708 3290
rect 11760 3238 11772 3290
rect 11824 3238 11836 3290
rect 11888 3238 11900 3290
rect 11952 3238 22338 3290
rect 22390 3238 22402 3290
rect 22454 3238 22466 3290
rect 22518 3238 22530 3290
rect 22582 3238 22594 3290
rect 22646 3238 33032 3290
rect 33084 3238 33096 3290
rect 33148 3238 33160 3290
rect 33212 3238 33224 3290
rect 33276 3238 33288 3290
rect 33340 3238 43726 3290
rect 43778 3238 43790 3290
rect 43842 3238 43854 3290
rect 43906 3238 43918 3290
rect 43970 3238 43982 3290
rect 44034 3238 44040 3290
rect 1104 3216 44040 3238
rect 9306 3136 9312 3188
rect 9364 3136 9370 3188
rect 13906 3136 13912 3188
rect 13964 3136 13970 3188
rect 14553 3179 14611 3185
rect 14553 3145 14565 3179
rect 14599 3145 14611 3179
rect 14553 3139 14611 3145
rect 14829 3179 14887 3185
rect 14829 3145 14841 3179
rect 14875 3176 14887 3179
rect 14875 3148 18736 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 14568 3108 14596 3139
rect 18046 3108 18052 3120
rect 14568 3080 18052 3108
rect 18046 3068 18052 3080
rect 18104 3068 18110 3120
rect 18708 3108 18736 3148
rect 19150 3136 19156 3188
rect 19208 3136 19214 3188
rect 19334 3136 19340 3188
rect 19392 3136 19398 3188
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20036 3148 20760 3176
rect 20036 3136 20042 3148
rect 18708 3080 19196 3108
rect 9122 3000 9128 3052
rect 9180 3000 9186 3052
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 13998 3040 14004 3052
rect 13771 3012 14004 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 14642 3000 14648 3052
rect 14700 3000 14706 3052
rect 14918 3000 14924 3052
rect 14976 3000 14982 3052
rect 15378 3000 15384 3052
rect 15436 3000 15442 3052
rect 15654 3000 15660 3052
rect 15712 3000 15718 3052
rect 15930 3000 15936 3052
rect 15988 3000 15994 3052
rect 16206 3000 16212 3052
rect 16264 3000 16270 3052
rect 16482 3000 16488 3052
rect 16540 3000 16546 3052
rect 16942 3000 16948 3052
rect 17000 3000 17006 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 14090 2972 14096 2984
rect 13872 2944 14096 2972
rect 13872 2932 13878 2944
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 17052 2972 17080 3003
rect 17494 3000 17500 3052
rect 17552 3000 17558 3052
rect 17770 3000 17776 3052
rect 17828 3000 17834 3052
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3009 17923 3043
rect 17865 3003 17923 3009
rect 16776 2944 17080 2972
rect 15010 2864 15016 2916
rect 15068 2904 15074 2916
rect 16776 2913 16804 2944
rect 16761 2907 16819 2913
rect 15068 2876 15240 2904
rect 15068 2864 15074 2876
rect 15102 2796 15108 2848
rect 15160 2796 15166 2848
rect 15212 2845 15240 2876
rect 16761 2873 16773 2907
rect 16807 2873 16819 2907
rect 17589 2907 17647 2913
rect 16761 2867 16819 2873
rect 17236 2876 17540 2904
rect 15197 2839 15255 2845
rect 15197 2805 15209 2839
rect 15243 2805 15255 2839
rect 15197 2799 15255 2805
rect 15286 2796 15292 2848
rect 15344 2836 15350 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15344 2808 15485 2836
rect 15344 2796 15350 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 15562 2796 15568 2848
rect 15620 2836 15626 2848
rect 15749 2839 15807 2845
rect 15749 2836 15761 2839
rect 15620 2808 15761 2836
rect 15620 2796 15626 2808
rect 15749 2805 15761 2808
rect 15795 2805 15807 2839
rect 15749 2799 15807 2805
rect 15838 2796 15844 2848
rect 15896 2836 15902 2848
rect 16025 2839 16083 2845
rect 16025 2836 16037 2839
rect 15896 2808 16037 2836
rect 15896 2796 15902 2808
rect 16025 2805 16037 2808
rect 16071 2805 16083 2839
rect 16025 2799 16083 2805
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 17236 2845 17264 2876
rect 17512 2848 17540 2876
rect 17589 2873 17601 2907
rect 17635 2904 17647 2907
rect 17880 2904 17908 3003
rect 18138 3000 18144 3052
rect 18196 3000 18202 3052
rect 18598 3000 18604 3052
rect 18656 3000 18662 3052
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3040 18751 3043
rect 18782 3040 18788 3052
rect 18739 3012 18788 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 18969 3043 19027 3049
rect 18969 3009 18981 3043
rect 19015 3009 19027 3043
rect 18969 3003 19027 3009
rect 18984 2972 19012 3003
rect 18432 2944 19012 2972
rect 19168 2972 19196 3080
rect 19245 3043 19303 3049
rect 19245 3009 19257 3043
rect 19291 3040 19303 3043
rect 19352 3040 19380 3136
rect 20732 3117 20760 3148
rect 20806 3136 20812 3188
rect 20864 3136 20870 3188
rect 21450 3136 21456 3188
rect 21508 3136 21514 3188
rect 22002 3136 22008 3188
rect 22060 3176 22066 3188
rect 22060 3148 22784 3176
rect 22060 3136 22066 3148
rect 20717 3111 20775 3117
rect 20717 3077 20729 3111
rect 20763 3077 20775 3111
rect 20824 3108 20852 3136
rect 21269 3111 21327 3117
rect 21269 3108 21281 3111
rect 20824 3080 21281 3108
rect 20717 3071 20775 3077
rect 21269 3077 21281 3080
rect 21315 3077 21327 3111
rect 21468 3108 21496 3136
rect 22756 3117 22784 3148
rect 22922 3136 22928 3188
rect 22980 3136 22986 3188
rect 24029 3179 24087 3185
rect 24029 3145 24041 3179
rect 24075 3176 24087 3179
rect 24075 3148 24716 3176
rect 24075 3145 24087 3148
rect 24029 3139 24087 3145
rect 22189 3111 22247 3117
rect 22189 3108 22201 3111
rect 21468 3080 22201 3108
rect 21269 3071 21327 3077
rect 22189 3077 22201 3080
rect 22235 3077 22247 3111
rect 22189 3071 22247 3077
rect 22741 3111 22799 3117
rect 22741 3077 22753 3111
rect 22787 3077 22799 3111
rect 22940 3108 22968 3136
rect 23293 3111 23351 3117
rect 23293 3108 23305 3111
rect 22940 3080 23305 3108
rect 22741 3071 22799 3077
rect 23293 3077 23305 3080
rect 23339 3077 23351 3111
rect 23293 3071 23351 3077
rect 24394 3068 24400 3120
rect 24452 3108 24458 3120
rect 24688 3117 24716 3148
rect 25222 3136 25228 3188
rect 25280 3136 25286 3188
rect 26326 3136 26332 3188
rect 26384 3176 26390 3188
rect 26384 3148 27660 3176
rect 26384 3136 26390 3148
rect 24673 3111 24731 3117
rect 24452 3080 24624 3108
rect 24452 3068 24458 3080
rect 19291 3012 19380 3040
rect 19291 3009 19303 3012
rect 19245 3003 19303 3009
rect 19610 3000 19616 3052
rect 19668 3000 19674 3052
rect 19886 3000 19892 3052
rect 19944 3040 19950 3052
rect 20165 3043 20223 3049
rect 20165 3040 20177 3043
rect 19944 3012 20177 3040
rect 19944 3000 19950 3012
rect 20165 3009 20177 3012
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 20806 3000 20812 3052
rect 20864 3040 20870 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 20864 3012 22017 3040
rect 20864 3000 20870 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 23750 3000 23756 3052
rect 23808 3040 23814 3052
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 23808 3012 23949 3040
rect 23808 3000 23814 3012
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 24210 3000 24216 3052
rect 24268 3000 24274 3052
rect 24486 3000 24492 3052
rect 24544 3000 24550 3052
rect 24596 3040 24624 3080
rect 24673 3077 24685 3111
rect 24719 3077 24731 3111
rect 25240 3108 25268 3136
rect 25240 3080 26372 3108
rect 24673 3071 24731 3077
rect 25225 3043 25283 3049
rect 25225 3040 25237 3043
rect 24596 3012 25237 3040
rect 25225 3009 25237 3012
rect 25271 3009 25283 3043
rect 25225 3003 25283 3009
rect 25777 3043 25835 3049
rect 25777 3009 25789 3043
rect 25823 3040 25835 3043
rect 26234 3040 26240 3052
rect 25823 3012 26240 3040
rect 25823 3009 25835 3012
rect 25777 3003 25835 3009
rect 26234 3000 26240 3012
rect 26292 3000 26298 3052
rect 26344 3049 26372 3080
rect 26694 3068 26700 3120
rect 26752 3068 26758 3120
rect 26878 3068 26884 3120
rect 26936 3108 26942 3120
rect 27632 3117 27660 3148
rect 28074 3136 28080 3188
rect 28132 3136 28138 3188
rect 28626 3136 28632 3188
rect 28684 3176 28690 3188
rect 28684 3148 29868 3176
rect 28684 3136 28690 3148
rect 27617 3111 27675 3117
rect 26936 3080 27568 3108
rect 26936 3068 26942 3080
rect 26329 3043 26387 3049
rect 26329 3009 26341 3043
rect 26375 3009 26387 3043
rect 26712 3040 26740 3068
rect 27065 3043 27123 3049
rect 27065 3040 27077 3043
rect 26712 3012 27077 3040
rect 26329 3003 26387 3009
rect 27065 3009 27077 3012
rect 27111 3009 27123 3043
rect 27540 3040 27568 3080
rect 27617 3077 27629 3111
rect 27663 3077 27675 3111
rect 28092 3108 28120 3136
rect 29840 3117 29868 3148
rect 30558 3136 30564 3188
rect 30616 3176 30622 3188
rect 31573 3179 31631 3185
rect 31573 3176 31585 3179
rect 30616 3148 31585 3176
rect 30616 3136 30622 3148
rect 31573 3145 31585 3148
rect 31619 3145 31631 3179
rect 31573 3139 31631 3145
rect 33042 3136 33048 3188
rect 33100 3176 33106 3188
rect 33965 3179 34023 3185
rect 33965 3176 33977 3179
rect 33100 3148 33977 3176
rect 33100 3136 33106 3148
rect 33965 3145 33977 3148
rect 34011 3145 34023 3179
rect 33965 3139 34023 3145
rect 34514 3136 34520 3188
rect 34572 3176 34578 3188
rect 35069 3179 35127 3185
rect 35069 3176 35081 3179
rect 34572 3148 35081 3176
rect 34572 3136 34578 3148
rect 35069 3145 35081 3148
rect 35115 3145 35127 3179
rect 35069 3139 35127 3145
rect 35437 3179 35495 3185
rect 35437 3145 35449 3179
rect 35483 3176 35495 3179
rect 35526 3176 35532 3188
rect 35483 3148 35532 3176
rect 35483 3145 35495 3148
rect 35437 3139 35495 3145
rect 35526 3136 35532 3148
rect 35584 3136 35590 3188
rect 35618 3136 35624 3188
rect 35676 3176 35682 3188
rect 38105 3179 38163 3185
rect 38105 3176 38117 3179
rect 35676 3148 38117 3176
rect 35676 3136 35682 3148
rect 38105 3145 38117 3148
rect 38151 3145 38163 3179
rect 38105 3139 38163 3145
rect 29273 3111 29331 3117
rect 29273 3108 29285 3111
rect 28092 3080 29285 3108
rect 27617 3071 27675 3077
rect 29273 3077 29285 3080
rect 29319 3077 29331 3111
rect 29273 3071 29331 3077
rect 29825 3111 29883 3117
rect 29825 3077 29837 3111
rect 29871 3077 29883 3111
rect 30929 3111 30987 3117
rect 30929 3108 30941 3111
rect 29825 3071 29883 3077
rect 29932 3080 30941 3108
rect 28169 3043 28227 3049
rect 28169 3040 28181 3043
rect 27540 3012 28181 3040
rect 27065 3003 27123 3009
rect 28169 3009 28181 3012
rect 28215 3009 28227 3043
rect 28169 3003 28227 3009
rect 28721 3043 28779 3049
rect 28721 3009 28733 3043
rect 28767 3040 28779 3043
rect 28902 3040 28908 3052
rect 28767 3012 28908 3040
rect 28767 3009 28779 3012
rect 28721 3003 28779 3009
rect 28902 3000 28908 3012
rect 28960 3000 28966 3052
rect 28994 3000 29000 3052
rect 29052 3040 29058 3052
rect 29932 3040 29960 3080
rect 30929 3077 30941 3080
rect 30975 3077 30987 3111
rect 30929 3071 30987 3077
rect 33410 3068 33416 3120
rect 33468 3108 33474 3120
rect 34425 3111 34483 3117
rect 34425 3108 34437 3111
rect 33468 3080 34437 3108
rect 33468 3068 33474 3080
rect 34425 3077 34437 3080
rect 34471 3077 34483 3111
rect 34425 3071 34483 3077
rect 34974 3068 34980 3120
rect 35032 3068 35038 3120
rect 35250 3068 35256 3120
rect 35308 3108 35314 3120
rect 35308 3080 36124 3108
rect 35308 3068 35314 3080
rect 29052 3012 29960 3040
rect 29052 3000 29058 3012
rect 30006 3000 30012 3052
rect 30064 3040 30070 3052
rect 30377 3043 30435 3049
rect 30377 3040 30389 3043
rect 30064 3012 30389 3040
rect 30064 3000 30070 3012
rect 30377 3009 30389 3012
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 31481 3043 31539 3049
rect 31481 3009 31493 3043
rect 31527 3009 31539 3043
rect 31481 3003 31539 3009
rect 19334 2972 19340 2984
rect 19168 2944 19340 2972
rect 17635 2876 17908 2904
rect 17635 2873 17647 2876
rect 17589 2867 17647 2873
rect 18322 2864 18328 2916
rect 18380 2864 18386 2916
rect 18432 2913 18460 2944
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 23566 2972 23572 2984
rect 19444 2944 23572 2972
rect 19444 2913 19472 2944
rect 23566 2932 23572 2944
rect 23624 2932 23630 2984
rect 24854 2972 24860 2984
rect 23768 2944 24860 2972
rect 18417 2907 18475 2913
rect 18417 2873 18429 2907
rect 18463 2873 18475 2907
rect 19429 2907 19487 2913
rect 18417 2867 18475 2873
rect 18800 2876 19288 2904
rect 16301 2839 16359 2845
rect 16301 2836 16313 2839
rect 16172 2808 16313 2836
rect 16172 2796 16178 2808
rect 16301 2805 16313 2808
rect 16347 2805 16359 2839
rect 16301 2799 16359 2805
rect 17221 2839 17279 2845
rect 17221 2805 17233 2839
rect 17267 2805 17279 2839
rect 17221 2799 17279 2805
rect 17310 2796 17316 2848
rect 17368 2796 17374 2848
rect 17494 2796 17500 2848
rect 17552 2796 17558 2848
rect 18049 2839 18107 2845
rect 18049 2805 18061 2839
rect 18095 2836 18107 2839
rect 18800 2836 18828 2876
rect 18095 2808 18828 2836
rect 18095 2805 18107 2808
rect 18049 2799 18107 2805
rect 18874 2796 18880 2848
rect 18932 2796 18938 2848
rect 19260 2836 19288 2876
rect 19429 2873 19441 2907
rect 19475 2873 19487 2907
rect 19429 2867 19487 2873
rect 19794 2864 19800 2916
rect 19852 2864 19858 2916
rect 20990 2904 20996 2916
rect 20180 2876 20996 2904
rect 20180 2836 20208 2876
rect 20990 2864 20996 2876
rect 21048 2864 21054 2916
rect 22002 2864 22008 2916
rect 22060 2904 22066 2916
rect 22060 2876 22324 2904
rect 22060 2864 22066 2876
rect 19260 2808 20208 2836
rect 20254 2796 20260 2848
rect 20312 2796 20318 2848
rect 20622 2796 20628 2848
rect 20680 2836 20686 2848
rect 20809 2839 20867 2845
rect 20809 2836 20821 2839
rect 20680 2808 20821 2836
rect 20680 2796 20686 2808
rect 20809 2805 20821 2808
rect 20855 2805 20867 2839
rect 20809 2799 20867 2805
rect 21358 2796 21364 2848
rect 21416 2796 21422 2848
rect 21821 2839 21879 2845
rect 21821 2805 21833 2839
rect 21867 2836 21879 2839
rect 22094 2836 22100 2848
rect 21867 2808 22100 2836
rect 21867 2805 21879 2808
rect 21821 2799 21879 2805
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 22296 2845 22324 2876
rect 22281 2839 22339 2845
rect 22281 2805 22293 2839
rect 22327 2805 22339 2839
rect 22281 2799 22339 2805
rect 22830 2796 22836 2848
rect 22888 2796 22894 2848
rect 23106 2796 23112 2848
rect 23164 2836 23170 2848
rect 23768 2845 23796 2944
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 31496 2972 31524 3003
rect 32306 3000 32312 3052
rect 32364 3040 32370 3052
rect 32769 3043 32827 3049
rect 32769 3040 32781 3043
rect 32364 3012 32781 3040
rect 32364 3000 32370 3012
rect 32769 3009 32781 3012
rect 32815 3009 32827 3043
rect 32769 3003 32827 3009
rect 33321 3043 33379 3049
rect 33321 3009 33333 3043
rect 33367 3040 33379 3043
rect 33686 3040 33692 3052
rect 33367 3012 33692 3040
rect 33367 3009 33379 3012
rect 33321 3003 33379 3009
rect 33686 3000 33692 3012
rect 33744 3000 33750 3052
rect 33778 3000 33784 3052
rect 33836 3040 33842 3052
rect 33873 3043 33931 3049
rect 33873 3040 33885 3043
rect 33836 3012 33885 3040
rect 33836 3000 33842 3012
rect 33873 3009 33885 3012
rect 33919 3009 33931 3043
rect 33873 3003 33931 3009
rect 35342 3000 35348 3052
rect 35400 3000 35406 3052
rect 36096 3049 36124 3080
rect 36814 3068 36820 3120
rect 36872 3068 36878 3120
rect 35805 3043 35863 3049
rect 35805 3040 35817 3043
rect 35452 3012 35817 3040
rect 29144 2944 31524 2972
rect 29144 2932 29150 2944
rect 34698 2932 34704 2984
rect 34756 2972 34762 2984
rect 35452 2972 35480 3012
rect 35805 3009 35817 3012
rect 35851 3009 35863 3043
rect 35805 3003 35863 3009
rect 36081 3043 36139 3049
rect 36081 3009 36093 3043
rect 36127 3009 36139 3043
rect 36081 3003 36139 3009
rect 36173 3043 36231 3049
rect 36173 3009 36185 3043
rect 36219 3009 36231 3043
rect 36173 3003 36231 3009
rect 34756 2944 35480 2972
rect 34756 2932 34762 2944
rect 35710 2932 35716 2984
rect 35768 2972 35774 2984
rect 36188 2972 36216 3003
rect 35768 2944 36216 2972
rect 35768 2932 35774 2944
rect 24946 2904 24952 2916
rect 24320 2876 24952 2904
rect 24320 2845 24348 2876
rect 24946 2864 24952 2876
rect 25004 2864 25010 2916
rect 26970 2864 26976 2916
rect 27028 2904 27034 2916
rect 27028 2876 27292 2904
rect 27028 2864 27034 2876
rect 23385 2839 23443 2845
rect 23385 2836 23397 2839
rect 23164 2808 23397 2836
rect 23164 2796 23170 2808
rect 23385 2805 23397 2808
rect 23431 2805 23443 2839
rect 23385 2799 23443 2805
rect 23753 2839 23811 2845
rect 23753 2805 23765 2839
rect 23799 2805 23811 2839
rect 23753 2799 23811 2805
rect 24305 2839 24363 2845
rect 24305 2805 24317 2839
rect 24351 2805 24363 2839
rect 24305 2799 24363 2805
rect 24486 2796 24492 2848
rect 24544 2836 24550 2848
rect 24765 2839 24823 2845
rect 24765 2836 24777 2839
rect 24544 2808 24777 2836
rect 24544 2796 24550 2808
rect 24765 2805 24777 2808
rect 24811 2805 24823 2839
rect 24765 2799 24823 2805
rect 25038 2796 25044 2848
rect 25096 2836 25102 2848
rect 25317 2839 25375 2845
rect 25317 2836 25329 2839
rect 25096 2808 25329 2836
rect 25096 2796 25102 2808
rect 25317 2805 25329 2808
rect 25363 2805 25375 2839
rect 25317 2799 25375 2805
rect 25590 2796 25596 2848
rect 25648 2836 25654 2848
rect 25869 2839 25927 2845
rect 25869 2836 25881 2839
rect 25648 2808 25881 2836
rect 25648 2796 25654 2808
rect 25869 2805 25881 2808
rect 25915 2805 25927 2839
rect 25869 2799 25927 2805
rect 26050 2796 26056 2848
rect 26108 2836 26114 2848
rect 26421 2839 26479 2845
rect 26421 2836 26433 2839
rect 26108 2808 26433 2836
rect 26108 2796 26114 2808
rect 26421 2805 26433 2808
rect 26467 2805 26479 2839
rect 26421 2799 26479 2805
rect 26602 2796 26608 2848
rect 26660 2836 26666 2848
rect 27157 2839 27215 2845
rect 27157 2836 27169 2839
rect 26660 2808 27169 2836
rect 26660 2796 26666 2808
rect 27157 2805 27169 2808
rect 27203 2805 27215 2839
rect 27264 2836 27292 2876
rect 27522 2864 27528 2916
rect 27580 2904 27586 2916
rect 27580 2876 28304 2904
rect 27580 2864 27586 2876
rect 28276 2845 28304 2876
rect 29730 2864 29736 2916
rect 29788 2904 29794 2916
rect 29788 2876 30052 2904
rect 29788 2864 29794 2876
rect 27709 2839 27767 2845
rect 27709 2836 27721 2839
rect 27264 2808 27721 2836
rect 27157 2799 27215 2805
rect 27709 2805 27721 2808
rect 27755 2805 27767 2839
rect 27709 2799 27767 2805
rect 28261 2839 28319 2845
rect 28261 2805 28273 2839
rect 28307 2805 28319 2839
rect 28261 2799 28319 2805
rect 28350 2796 28356 2848
rect 28408 2836 28414 2848
rect 28813 2839 28871 2845
rect 28813 2836 28825 2839
rect 28408 2808 28825 2836
rect 28408 2796 28414 2808
rect 28813 2805 28825 2808
rect 28859 2805 28871 2839
rect 28813 2799 28871 2805
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 29365 2839 29423 2845
rect 29365 2836 29377 2839
rect 28960 2808 29377 2836
rect 28960 2796 28966 2808
rect 29365 2805 29377 2808
rect 29411 2805 29423 2839
rect 29365 2799 29423 2805
rect 29454 2796 29460 2848
rect 29512 2836 29518 2848
rect 29917 2839 29975 2845
rect 29917 2836 29929 2839
rect 29512 2808 29929 2836
rect 29512 2796 29518 2808
rect 29917 2805 29929 2808
rect 29963 2805 29975 2839
rect 30024 2836 30052 2876
rect 30282 2864 30288 2916
rect 30340 2904 30346 2916
rect 30340 2876 31064 2904
rect 30340 2864 30346 2876
rect 31036 2845 31064 2876
rect 31938 2864 31944 2916
rect 31996 2904 32002 2916
rect 31996 2876 32444 2904
rect 31996 2864 32002 2876
rect 30469 2839 30527 2845
rect 30469 2836 30481 2839
rect 30024 2808 30481 2836
rect 29917 2799 29975 2805
rect 30469 2805 30481 2808
rect 30515 2805 30527 2839
rect 30469 2799 30527 2805
rect 31021 2839 31079 2845
rect 31021 2805 31033 2839
rect 31067 2805 31079 2839
rect 31021 2799 31079 2805
rect 32306 2796 32312 2848
rect 32364 2796 32370 2848
rect 32416 2836 32444 2876
rect 32490 2864 32496 2916
rect 32548 2904 32554 2916
rect 32548 2876 33456 2904
rect 32548 2864 32554 2876
rect 33428 2845 33456 2876
rect 33594 2864 33600 2916
rect 33652 2904 33658 2916
rect 35621 2907 35679 2913
rect 33652 2876 34560 2904
rect 33652 2864 33658 2876
rect 34532 2845 34560 2876
rect 35621 2873 35633 2907
rect 35667 2904 35679 2907
rect 35986 2904 35992 2916
rect 35667 2876 35992 2904
rect 35667 2873 35679 2876
rect 35621 2867 35679 2873
rect 35986 2864 35992 2876
rect 36044 2864 36050 2916
rect 36832 2904 36860 3068
rect 37734 3000 37740 3052
rect 37792 3040 37798 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37792 3012 38025 3040
rect 37792 3000 37798 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 38289 3043 38347 3049
rect 38289 3009 38301 3043
rect 38335 3009 38347 3043
rect 38289 3003 38347 3009
rect 38304 2972 38332 3003
rect 38838 3000 38844 3052
rect 38896 3040 38902 3052
rect 39117 3043 39175 3049
rect 39117 3040 39129 3043
rect 38896 3012 39129 3040
rect 38896 3000 38902 3012
rect 39117 3009 39129 3012
rect 39163 3009 39175 3043
rect 39117 3003 39175 3009
rect 39390 3000 39396 3052
rect 39448 3000 39454 3052
rect 40126 2972 40132 2984
rect 38304 2944 40132 2972
rect 40126 2932 40132 2944
rect 40184 2932 40190 2984
rect 37829 2907 37887 2913
rect 37829 2904 37841 2907
rect 36832 2876 37841 2904
rect 37829 2873 37841 2876
rect 37875 2873 37887 2907
rect 37829 2867 37887 2873
rect 32861 2839 32919 2845
rect 32861 2836 32873 2839
rect 32416 2808 32873 2836
rect 32861 2805 32873 2808
rect 32907 2805 32919 2839
rect 32861 2799 32919 2805
rect 33413 2839 33471 2845
rect 33413 2805 33425 2839
rect 33459 2805 33471 2839
rect 33413 2799 33471 2805
rect 34517 2839 34575 2845
rect 34517 2805 34529 2839
rect 34563 2805 34575 2839
rect 34517 2799 34575 2805
rect 35897 2839 35955 2845
rect 35897 2805 35909 2839
rect 35943 2836 35955 2839
rect 36078 2836 36084 2848
rect 35943 2808 36084 2836
rect 35943 2805 35955 2808
rect 35897 2799 35955 2805
rect 36078 2796 36084 2808
rect 36136 2796 36142 2848
rect 36354 2796 36360 2848
rect 36412 2796 36418 2848
rect 37182 2796 37188 2848
rect 37240 2836 37246 2848
rect 38746 2836 38752 2848
rect 37240 2808 38752 2836
rect 37240 2796 37246 2808
rect 38746 2796 38752 2808
rect 38804 2796 38810 2848
rect 38933 2839 38991 2845
rect 38933 2805 38945 2839
rect 38979 2836 38991 2839
rect 39114 2836 39120 2848
rect 38979 2808 39120 2836
rect 38979 2805 38991 2808
rect 38933 2799 38991 2805
rect 39114 2796 39120 2808
rect 39172 2796 39178 2848
rect 39209 2839 39267 2845
rect 39209 2805 39221 2839
rect 39255 2836 39267 2839
rect 40402 2836 40408 2848
rect 39255 2808 40408 2836
rect 39255 2805 39267 2808
rect 39209 2799 39267 2805
rect 40402 2796 40408 2808
rect 40460 2796 40466 2848
rect 1104 2746 43884 2768
rect 1104 2694 6297 2746
rect 6349 2694 6361 2746
rect 6413 2694 6425 2746
rect 6477 2694 6489 2746
rect 6541 2694 6553 2746
rect 6605 2694 16991 2746
rect 17043 2694 17055 2746
rect 17107 2694 17119 2746
rect 17171 2694 17183 2746
rect 17235 2694 17247 2746
rect 17299 2694 27685 2746
rect 27737 2694 27749 2746
rect 27801 2694 27813 2746
rect 27865 2694 27877 2746
rect 27929 2694 27941 2746
rect 27993 2694 38379 2746
rect 38431 2694 38443 2746
rect 38495 2694 38507 2746
rect 38559 2694 38571 2746
rect 38623 2694 38635 2746
rect 38687 2694 43884 2746
rect 1104 2672 43884 2694
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 5675 2604 6316 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 4801 2567 4859 2573
rect 4801 2533 4813 2567
rect 4847 2564 4859 2567
rect 5902 2564 5908 2576
rect 4847 2536 5908 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 6178 2524 6184 2576
rect 6236 2524 6242 2576
rect 6288 2564 6316 2604
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 8662 2632 8668 2644
rect 6604 2604 8668 2632
rect 6604 2592 6610 2604
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 8757 2635 8815 2641
rect 8757 2601 8769 2635
rect 8803 2601 8815 2635
rect 9214 2632 9220 2644
rect 8757 2595 8815 2601
rect 9048 2604 9220 2632
rect 7101 2567 7159 2573
rect 6288 2536 6914 2564
rect 5534 2496 5540 2508
rect 5184 2468 5540 2496
rect 5184 2437 5212 2468
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5810 2496 5816 2508
rect 5644 2468 5816 2496
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5169 2431 5227 2437
rect 4939 2400 5120 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 4632 2360 4660 2391
rect 4982 2360 4988 2372
rect 4632 2332 4988 2360
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 5092 2360 5120 2400
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5644 2428 5672 2468
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 6270 2456 6276 2508
rect 6328 2456 6334 2508
rect 6730 2496 6736 2508
rect 6380 2468 6736 2496
rect 5491 2400 5672 2428
rect 5721 2431 5779 2437
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5721 2397 5733 2431
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6288 2428 6316 2456
rect 6380 2437 6408 2468
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 6886 2496 6914 2536
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 8294 2564 8300 2576
rect 7147 2536 8300 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 8772 2508 8800 2595
rect 9048 2564 9076 2604
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9398 2592 9404 2644
rect 9456 2592 9462 2644
rect 9950 2592 9956 2644
rect 10008 2592 10014 2644
rect 10226 2592 10232 2644
rect 10284 2592 10290 2644
rect 11054 2592 11060 2644
rect 11112 2592 11118 2644
rect 13262 2632 13268 2644
rect 11716 2604 13268 2632
rect 11716 2573 11744 2604
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13814 2632 13820 2644
rect 13372 2604 13820 2632
rect 9125 2567 9183 2573
rect 9125 2564 9137 2567
rect 9048 2536 9137 2564
rect 9125 2533 9137 2536
rect 9171 2533 9183 2567
rect 9125 2527 9183 2533
rect 9493 2567 9551 2573
rect 9493 2533 9505 2567
rect 9539 2564 9551 2567
rect 11701 2567 11759 2573
rect 9539 2536 11468 2564
rect 9539 2533 9551 2536
rect 9493 2527 9551 2533
rect 6886 2468 8248 2496
rect 8220 2440 8248 2468
rect 8754 2456 8760 2508
rect 8812 2456 8818 2508
rect 9858 2496 9864 2508
rect 9232 2468 9864 2496
rect 6043 2400 6316 2428
rect 6365 2431 6423 2437
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 5258 2360 5264 2372
rect 5092 2332 5264 2360
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 4890 2252 4896 2304
rect 4948 2292 4954 2304
rect 5077 2295 5135 2301
rect 5077 2292 5089 2295
rect 4948 2264 5089 2292
rect 4948 2252 4954 2264
rect 5077 2261 5089 2264
rect 5123 2261 5135 2295
rect 5077 2255 5135 2261
rect 5353 2295 5411 2301
rect 5353 2261 5365 2295
rect 5399 2292 5411 2295
rect 5534 2292 5540 2304
rect 5399 2264 5540 2292
rect 5399 2261 5411 2264
rect 5353 2255 5411 2261
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 5626 2252 5632 2304
rect 5684 2292 5690 2304
rect 5736 2292 5764 2391
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2397 6699 2431
rect 6641 2391 6699 2397
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7193 2431 7251 2437
rect 6963 2400 7144 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 6564 2360 6592 2388
rect 6380 2332 6592 2360
rect 6656 2360 6684 2391
rect 7006 2360 7012 2372
rect 6656 2332 7012 2360
rect 5684 2264 5764 2292
rect 5905 2295 5963 2301
rect 5684 2252 5690 2264
rect 5905 2261 5917 2295
rect 5951 2292 5963 2295
rect 6380 2292 6408 2332
rect 7006 2320 7012 2332
rect 7064 2320 7070 2372
rect 7116 2360 7144 2400
rect 7193 2397 7205 2431
rect 7239 2428 7251 2431
rect 7374 2428 7380 2440
rect 7239 2400 7380 2428
rect 7239 2397 7251 2400
rect 7193 2391 7251 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7650 2428 7656 2440
rect 7515 2400 7656 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 7926 2428 7932 2440
rect 7791 2400 7932 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 7282 2360 7288 2372
rect 7116 2332 7288 2360
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 7834 2360 7840 2372
rect 7668 2332 7840 2360
rect 5951 2264 6408 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 6546 2252 6552 2304
rect 6604 2252 6610 2304
rect 6822 2252 6828 2304
rect 6880 2252 6886 2304
rect 7374 2252 7380 2304
rect 7432 2252 7438 2304
rect 7668 2301 7696 2332
rect 7834 2320 7840 2332
rect 7892 2320 7898 2372
rect 8036 2360 8064 2391
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2428 8355 2431
rect 8343 2400 8524 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 8386 2360 8392 2372
rect 8036 2332 8392 2360
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 8496 2360 8524 2400
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 9232 2437 9260 2468
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 10410 2496 10416 2508
rect 9968 2468 10416 2496
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 9968 2428 9996 2468
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 10962 2496 10968 2508
rect 10520 2468 10968 2496
rect 9815 2400 9996 2428
rect 10045 2431 10103 2437
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10321 2431 10379 2437
rect 10091 2400 10272 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 8662 2360 8668 2372
rect 8496 2332 8668 2360
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 8956 2360 8984 2391
rect 9582 2360 9588 2372
rect 8956 2332 9588 2360
rect 9582 2320 9588 2332
rect 9640 2320 9646 2372
rect 9692 2360 9720 2391
rect 10134 2360 10140 2372
rect 9692 2332 10140 2360
rect 10134 2320 10140 2332
rect 10192 2320 10198 2372
rect 10244 2360 10272 2400
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10520 2428 10548 2468
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 11440 2440 11468 2536
rect 11701 2533 11713 2567
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 11974 2524 11980 2576
rect 12032 2524 12038 2576
rect 12250 2524 12256 2576
rect 12308 2524 12314 2576
rect 12526 2524 12532 2576
rect 12584 2524 12590 2576
rect 13081 2567 13139 2573
rect 13081 2533 13093 2567
rect 13127 2564 13139 2567
rect 13372 2564 13400 2604
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 13906 2592 13912 2644
rect 13964 2592 13970 2644
rect 14093 2635 14151 2641
rect 14093 2601 14105 2635
rect 14139 2632 14151 2635
rect 14182 2632 14188 2644
rect 14139 2604 14188 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 18138 2632 18144 2644
rect 17267 2604 18144 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19610 2632 19616 2644
rect 18800 2604 19616 2632
rect 13127 2536 13400 2564
rect 13449 2567 13507 2573
rect 13127 2533 13139 2536
rect 13081 2527 13139 2533
rect 13449 2533 13461 2567
rect 13495 2564 13507 2567
rect 16942 2564 16948 2576
rect 13495 2536 13768 2564
rect 13495 2533 13507 2536
rect 13449 2527 13507 2533
rect 12802 2496 12808 2508
rect 12360 2468 12808 2496
rect 10367 2400 10548 2428
rect 10597 2431 10655 2437
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 10873 2431 10931 2437
rect 10643 2400 10824 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 10686 2360 10692 2372
rect 10244 2332 10692 2360
rect 10686 2320 10692 2332
rect 10744 2320 10750 2372
rect 10796 2360 10824 2400
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 11054 2428 11060 2440
rect 10919 2400 11060 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11422 2388 11428 2440
rect 11480 2388 11486 2440
rect 12360 2437 12388 2468
rect 12802 2456 12808 2468
rect 12860 2456 12866 2508
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 11793 2431 11851 2437
rect 11793 2397 11805 2431
rect 11839 2428 11851 2431
rect 12069 2431 12127 2437
rect 11839 2400 12020 2428
rect 11839 2397 11851 2400
rect 11793 2391 11851 2397
rect 11238 2360 11244 2372
rect 10796 2332 11244 2360
rect 11238 2320 11244 2332
rect 11296 2320 11302 2372
rect 11532 2360 11560 2391
rect 11882 2360 11888 2372
rect 11532 2332 11888 2360
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 7653 2295 7711 2301
rect 7653 2261 7665 2295
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 7926 2252 7932 2304
rect 7984 2252 7990 2304
rect 8110 2252 8116 2304
rect 8168 2292 8174 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 8168 2264 8217 2292
rect 8168 2252 8174 2264
rect 8205 2261 8217 2264
rect 8251 2261 8263 2295
rect 8205 2255 8263 2261
rect 8481 2295 8539 2301
rect 8481 2261 8493 2295
rect 8527 2292 8539 2295
rect 10318 2292 10324 2304
rect 8527 2264 10324 2292
rect 8527 2261 8539 2264
rect 8481 2255 8539 2261
rect 10318 2252 10324 2264
rect 10376 2252 10382 2304
rect 10502 2252 10508 2304
rect 10560 2252 10566 2304
rect 10778 2252 10784 2304
rect 10836 2252 10842 2304
rect 11330 2252 11336 2304
rect 11388 2252 11394 2304
rect 11992 2292 12020 2400
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12345 2431 12403 2437
rect 12115 2400 12296 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12268 2360 12296 2400
rect 12345 2397 12357 2431
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2428 12679 2431
rect 12710 2428 12716 2440
rect 12667 2400 12716 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 13538 2428 13544 2440
rect 13219 2400 13544 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 12434 2360 12440 2372
rect 12268 2332 12440 2360
rect 12434 2320 12440 2332
rect 12492 2320 12498 2372
rect 12912 2360 12940 2391
rect 13538 2388 13544 2400
rect 13596 2388 13602 2440
rect 13740 2437 13768 2536
rect 13832 2536 16948 2564
rect 13832 2440 13860 2536
rect 16942 2524 16948 2536
rect 17000 2524 17006 2576
rect 17034 2524 17040 2576
rect 17092 2524 17098 2576
rect 17129 2567 17187 2573
rect 17129 2533 17141 2567
rect 17175 2564 17187 2567
rect 18049 2567 18107 2573
rect 17175 2536 18000 2564
rect 17175 2533 17187 2536
rect 17129 2527 17187 2533
rect 17052 2496 17080 2524
rect 17972 2496 18000 2536
rect 18049 2533 18061 2567
rect 18095 2564 18107 2567
rect 18800 2564 18828 2604
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 23658 2632 23664 2644
rect 19720 2604 23664 2632
rect 18095 2536 18828 2564
rect 19245 2567 19303 2573
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 19245 2533 19257 2567
rect 19291 2533 19303 2567
rect 19245 2527 19303 2533
rect 19150 2496 19156 2508
rect 15396 2468 17080 2496
rect 17420 2468 17908 2496
rect 17972 2468 19156 2496
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 13446 2360 13452 2372
rect 12912 2332 13452 2360
rect 13446 2320 13452 2332
rect 13504 2320 13510 2372
rect 13648 2360 13676 2391
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2428 14335 2431
rect 14826 2428 14832 2440
rect 14323 2400 14832 2428
rect 14323 2397 14335 2400
rect 14277 2391 14335 2397
rect 14826 2388 14832 2400
rect 14884 2388 14890 2440
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15010 2428 15016 2440
rect 14967 2400 15016 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15286 2428 15292 2440
rect 15243 2400 15292 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 15396 2360 15424 2468
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2428 15531 2431
rect 15562 2428 15568 2440
rect 15519 2400 15568 2428
rect 15519 2397 15531 2400
rect 15473 2391 15531 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2428 15807 2431
rect 15838 2428 15844 2440
rect 15795 2400 15844 2428
rect 15795 2397 15807 2400
rect 15749 2391 15807 2397
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2428 16083 2431
rect 16114 2428 16120 2440
rect 16071 2400 16120 2428
rect 16071 2397 16083 2400
rect 16025 2391 16083 2397
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 16298 2388 16304 2440
rect 16356 2388 16362 2440
rect 16666 2388 16672 2440
rect 16724 2388 16730 2440
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17310 2428 17316 2440
rect 16991 2400 17316 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 17420 2437 17448 2468
rect 17405 2431 17463 2437
rect 17405 2397 17417 2431
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 17678 2388 17684 2440
rect 17736 2388 17742 2440
rect 17770 2388 17776 2440
rect 17828 2388 17834 2440
rect 17880 2428 17908 2468
rect 19150 2456 19156 2468
rect 19208 2456 19214 2508
rect 19260 2496 19288 2527
rect 19334 2524 19340 2576
rect 19392 2564 19398 2576
rect 19720 2564 19748 2604
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 24762 2592 24768 2644
rect 24820 2632 24826 2644
rect 25685 2635 25743 2641
rect 25685 2632 25697 2635
rect 24820 2604 25697 2632
rect 24820 2592 24826 2604
rect 25685 2601 25697 2604
rect 25731 2601 25743 2635
rect 25685 2595 25743 2601
rect 26234 2592 26240 2644
rect 26292 2632 26298 2644
rect 26605 2635 26663 2641
rect 26605 2632 26617 2635
rect 26292 2604 26617 2632
rect 26292 2592 26298 2604
rect 26605 2601 26617 2604
rect 26651 2601 26663 2635
rect 26605 2595 26663 2601
rect 26878 2592 26884 2644
rect 26936 2632 26942 2644
rect 27709 2635 27767 2641
rect 27709 2632 27721 2635
rect 26936 2604 27721 2632
rect 26936 2592 26942 2604
rect 27709 2601 27721 2604
rect 27755 2601 27767 2635
rect 27709 2595 27767 2601
rect 28166 2592 28172 2644
rect 28224 2632 28230 2644
rect 28813 2635 28871 2641
rect 28813 2632 28825 2635
rect 28224 2604 28825 2632
rect 28224 2592 28230 2604
rect 28813 2601 28825 2604
rect 28859 2601 28871 2635
rect 28813 2595 28871 2601
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 29181 2635 29239 2641
rect 29181 2632 29193 2635
rect 29052 2604 29193 2632
rect 29052 2592 29058 2604
rect 29181 2601 29193 2604
rect 29227 2601 29239 2635
rect 29181 2595 29239 2601
rect 29638 2592 29644 2644
rect 29696 2632 29702 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 29696 2604 30849 2632
rect 29696 2592 29702 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 31754 2592 31760 2644
rect 31812 2592 31818 2644
rect 32861 2635 32919 2641
rect 32861 2601 32873 2635
rect 32907 2601 32919 2635
rect 32861 2595 32919 2601
rect 19392 2536 19748 2564
rect 21821 2567 21879 2573
rect 19392 2524 19398 2536
rect 21821 2533 21833 2567
rect 21867 2564 21879 2567
rect 21867 2536 23336 2564
rect 21867 2533 21879 2536
rect 21821 2527 21879 2533
rect 19260 2468 20208 2496
rect 17954 2428 17960 2440
rect 17880 2400 17960 2428
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18230 2388 18236 2440
rect 18288 2388 18294 2440
rect 18322 2388 18328 2440
rect 18380 2428 18386 2440
rect 18509 2431 18567 2437
rect 18509 2428 18521 2431
rect 18380 2400 18521 2428
rect 18380 2388 18386 2400
rect 18509 2397 18521 2400
rect 18555 2397 18567 2431
rect 18509 2391 18567 2397
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 19702 2428 19708 2440
rect 19659 2400 19708 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 19702 2388 19708 2400
rect 19760 2388 19766 2440
rect 19886 2388 19892 2440
rect 19944 2388 19950 2440
rect 20180 2437 20208 2468
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22336 2468 22784 2496
rect 22336 2456 22342 2468
rect 20165 2431 20223 2437
rect 20165 2397 20177 2431
rect 20211 2397 20223 2431
rect 20165 2391 20223 2397
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 20898 2428 20904 2440
rect 20763 2400 20904 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 20898 2388 20904 2400
rect 20956 2388 20962 2440
rect 21174 2388 21180 2440
rect 21232 2428 21238 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 21232 2400 21281 2428
rect 21232 2388 21238 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 21542 2388 21548 2440
rect 21600 2428 21606 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21600 2400 22017 2428
rect 21600 2388 21606 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 22370 2428 22376 2440
rect 22235 2400 22376 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 22370 2388 22376 2400
rect 22428 2388 22434 2440
rect 22756 2437 22784 2468
rect 23308 2437 23336 2536
rect 23566 2524 23572 2576
rect 23624 2524 23630 2576
rect 27430 2524 27436 2576
rect 27488 2564 27494 2576
rect 28353 2567 28411 2573
rect 28353 2564 28365 2567
rect 27488 2536 28365 2564
rect 27488 2524 27494 2536
rect 28353 2533 28365 2536
rect 28399 2533 28411 2567
rect 28353 2527 28411 2533
rect 28902 2524 28908 2576
rect 28960 2564 28966 2576
rect 30377 2567 30435 2573
rect 30377 2564 30389 2567
rect 28960 2536 30389 2564
rect 28960 2524 28966 2536
rect 30377 2533 30389 2536
rect 30423 2533 30435 2567
rect 30377 2527 30435 2533
rect 30926 2524 30932 2576
rect 30984 2564 30990 2576
rect 32876 2564 32904 2595
rect 33502 2592 33508 2644
rect 33560 2632 33566 2644
rect 34333 2635 34391 2641
rect 34333 2632 34345 2635
rect 33560 2604 34345 2632
rect 33560 2592 33566 2604
rect 34333 2601 34345 2604
rect 34379 2601 34391 2635
rect 34333 2595 34391 2601
rect 35342 2592 35348 2644
rect 35400 2632 35406 2644
rect 35400 2604 36584 2632
rect 35400 2592 35406 2604
rect 30984 2536 32904 2564
rect 30984 2524 30990 2536
rect 33410 2524 33416 2576
rect 33468 2564 33474 2576
rect 35529 2567 35587 2573
rect 35529 2564 35541 2567
rect 33468 2536 35541 2564
rect 33468 2524 33474 2536
rect 35529 2533 35541 2536
rect 35575 2533 35587 2567
rect 35529 2527 35587 2533
rect 35802 2524 35808 2576
rect 35860 2564 35866 2576
rect 36081 2567 36139 2573
rect 36081 2564 36093 2567
rect 35860 2536 36093 2564
rect 35860 2524 35866 2536
rect 36081 2533 36093 2536
rect 36127 2533 36139 2567
rect 36556 2564 36584 2604
rect 36722 2592 36728 2644
rect 36780 2592 36786 2644
rect 36817 2635 36875 2641
rect 36817 2601 36829 2635
rect 36863 2632 36875 2635
rect 36906 2632 36912 2644
rect 36863 2604 36912 2632
rect 36863 2601 36875 2604
rect 36817 2595 36875 2601
rect 36906 2592 36912 2604
rect 36964 2592 36970 2644
rect 36998 2592 37004 2644
rect 37056 2632 37062 2644
rect 39209 2635 39267 2641
rect 37056 2604 39160 2632
rect 37056 2592 37062 2604
rect 37277 2567 37335 2573
rect 37277 2564 37289 2567
rect 36556 2536 37289 2564
rect 36081 2527 36139 2533
rect 37277 2533 37289 2536
rect 37323 2533 37335 2567
rect 37277 2527 37335 2533
rect 37642 2524 37648 2576
rect 37700 2564 37706 2576
rect 39132 2573 39160 2604
rect 39209 2601 39221 2635
rect 39255 2632 39267 2635
rect 40034 2632 40040 2644
rect 39255 2604 40040 2632
rect 39255 2601 39267 2604
rect 39209 2595 39267 2601
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 40126 2592 40132 2644
rect 40184 2592 40190 2644
rect 40218 2592 40224 2644
rect 40276 2632 40282 2644
rect 40405 2635 40463 2641
rect 40405 2632 40417 2635
rect 40276 2604 40417 2632
rect 40276 2592 40282 2604
rect 40405 2601 40417 2604
rect 40451 2601 40463 2635
rect 40405 2595 40463 2601
rect 40494 2592 40500 2644
rect 40552 2592 40558 2644
rect 41233 2635 41291 2641
rect 41233 2601 41245 2635
rect 41279 2632 41291 2635
rect 41690 2632 41696 2644
rect 41279 2604 41696 2632
rect 41279 2601 41291 2604
rect 41233 2595 41291 2601
rect 41690 2592 41696 2604
rect 41748 2592 41754 2644
rect 42797 2635 42855 2641
rect 42797 2601 42809 2635
rect 42843 2632 42855 2635
rect 43162 2632 43168 2644
rect 42843 2604 43168 2632
rect 42843 2601 42855 2604
rect 42797 2595 42855 2601
rect 43162 2592 43168 2604
rect 43220 2592 43226 2644
rect 39117 2567 39175 2573
rect 37700 2536 38976 2564
rect 37700 2524 37706 2536
rect 23584 2496 23612 2524
rect 33597 2499 33655 2505
rect 33597 2496 33609 2499
rect 23584 2468 27660 2496
rect 22741 2431 22799 2437
rect 22741 2397 22753 2431
rect 22787 2397 22799 2431
rect 22741 2391 22799 2397
rect 23293 2431 23351 2437
rect 23293 2397 23305 2431
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23532 2400 23857 2428
rect 23532 2388 23538 2400
rect 23845 2397 23857 2400
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 23934 2388 23940 2440
rect 23992 2428 23998 2440
rect 24489 2431 24547 2437
rect 24489 2428 24501 2431
rect 23992 2400 24501 2428
rect 23992 2388 23998 2400
rect 24489 2397 24501 2400
rect 24535 2397 24547 2431
rect 24489 2391 24547 2397
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25041 2431 25099 2437
rect 25041 2428 25053 2431
rect 24912 2400 25053 2428
rect 24912 2388 24918 2400
rect 25041 2397 25053 2400
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 25682 2388 25688 2440
rect 25740 2428 25746 2440
rect 26145 2431 26203 2437
rect 26145 2428 26157 2431
rect 25740 2400 26157 2428
rect 25740 2388 25746 2400
rect 26145 2397 26157 2400
rect 26191 2397 26203 2431
rect 26145 2391 26203 2397
rect 26234 2388 26240 2440
rect 26292 2388 26298 2440
rect 26786 2388 26792 2440
rect 26844 2388 26850 2440
rect 27062 2388 27068 2440
rect 27120 2388 27126 2440
rect 27632 2428 27660 2468
rect 27908 2468 31340 2496
rect 27908 2440 27936 2468
rect 27632 2400 27844 2428
rect 16574 2360 16580 2372
rect 13648 2332 15056 2360
rect 15028 2304 15056 2332
rect 15212 2332 15424 2360
rect 16224 2332 16580 2360
rect 15212 2304 15240 2332
rect 12342 2292 12348 2304
rect 11992 2264 12348 2292
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 12802 2252 12808 2304
rect 12860 2252 12866 2304
rect 13357 2295 13415 2301
rect 13357 2261 13369 2295
rect 13403 2292 13415 2295
rect 14458 2292 14464 2304
rect 13403 2264 14464 2292
rect 13403 2261 13415 2264
rect 13357 2255 13415 2261
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14645 2295 14703 2301
rect 14645 2261 14657 2295
rect 14691 2292 14703 2295
rect 14826 2292 14832 2304
rect 14691 2264 14832 2292
rect 14691 2261 14703 2264
rect 14645 2255 14703 2261
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 15010 2252 15016 2304
rect 15068 2252 15074 2304
rect 15102 2252 15108 2304
rect 15160 2252 15166 2304
rect 15194 2252 15200 2304
rect 15252 2252 15258 2304
rect 15381 2295 15439 2301
rect 15381 2261 15393 2295
rect 15427 2292 15439 2295
rect 15562 2292 15568 2304
rect 15427 2264 15568 2292
rect 15427 2261 15439 2264
rect 15381 2255 15439 2261
rect 15562 2252 15568 2264
rect 15620 2252 15626 2304
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 15838 2292 15844 2304
rect 15703 2264 15844 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 15933 2295 15991 2301
rect 15933 2261 15945 2295
rect 15979 2292 15991 2295
rect 16114 2292 16120 2304
rect 15979 2264 16120 2292
rect 15979 2261 15991 2264
rect 15933 2255 15991 2261
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 16224 2301 16252 2332
rect 16574 2320 16580 2332
rect 16632 2320 16638 2372
rect 18693 2363 18751 2369
rect 18693 2360 18705 2363
rect 17512 2332 18705 2360
rect 16209 2295 16267 2301
rect 16209 2261 16221 2295
rect 16255 2261 16267 2295
rect 16209 2255 16267 2261
rect 16485 2295 16543 2301
rect 16485 2261 16497 2295
rect 16531 2292 16543 2295
rect 16666 2292 16672 2304
rect 16531 2264 16672 2292
rect 16531 2261 16543 2264
rect 16485 2255 16543 2261
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 17310 2292 17316 2304
rect 16899 2264 17316 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 17512 2301 17540 2332
rect 18693 2329 18705 2332
rect 18739 2329 18751 2363
rect 18693 2323 18751 2329
rect 19061 2363 19119 2369
rect 19061 2329 19073 2363
rect 19107 2360 19119 2363
rect 19518 2360 19524 2372
rect 19107 2332 19524 2360
rect 19107 2329 19119 2332
rect 19061 2323 19119 2329
rect 19518 2320 19524 2332
rect 19576 2320 19582 2372
rect 17497 2295 17555 2301
rect 17497 2261 17509 2295
rect 17543 2261 17555 2295
rect 17497 2255 17555 2261
rect 17957 2295 18015 2301
rect 17957 2261 17969 2295
rect 18003 2292 18015 2295
rect 18138 2292 18144 2304
rect 18003 2264 18144 2292
rect 18003 2261 18015 2264
rect 17957 2255 18015 2261
rect 18138 2252 18144 2264
rect 18196 2252 18202 2304
rect 18325 2295 18383 2301
rect 18325 2261 18337 2295
rect 18371 2292 18383 2295
rect 19904 2292 19932 2388
rect 19981 2363 20039 2369
rect 19981 2329 19993 2363
rect 20027 2360 20039 2363
rect 20346 2360 20352 2372
rect 20027 2332 20352 2360
rect 20027 2329 20039 2332
rect 19981 2323 20039 2329
rect 20346 2320 20352 2332
rect 20404 2320 20410 2372
rect 20533 2363 20591 2369
rect 20533 2329 20545 2363
rect 20579 2329 20591 2363
rect 20533 2323 20591 2329
rect 21085 2363 21143 2369
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21450 2360 21456 2372
rect 21131 2332 21456 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 18371 2264 19932 2292
rect 20548 2292 20576 2323
rect 21450 2320 21456 2332
rect 21508 2320 21514 2372
rect 21634 2320 21640 2372
rect 21692 2320 21698 2372
rect 24394 2320 24400 2372
rect 24452 2360 24458 2372
rect 24452 2332 24900 2360
rect 24452 2320 24458 2332
rect 20714 2292 20720 2304
rect 20548 2264 20720 2292
rect 18371 2261 18383 2264
rect 18325 2255 18383 2261
rect 20714 2252 20720 2264
rect 20772 2252 20778 2304
rect 22278 2252 22284 2304
rect 22336 2252 22342 2304
rect 22830 2252 22836 2304
rect 22888 2252 22894 2304
rect 23566 2252 23572 2304
rect 23624 2252 23630 2304
rect 23658 2252 23664 2304
rect 23716 2292 23722 2304
rect 23937 2295 23995 2301
rect 23937 2292 23949 2295
rect 23716 2264 23949 2292
rect 23716 2252 23722 2264
rect 23937 2261 23949 2264
rect 23983 2261 23995 2295
rect 23937 2255 23995 2261
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24084 2264 24593 2292
rect 24084 2252 24090 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24872 2292 24900 2332
rect 24946 2320 24952 2372
rect 25004 2360 25010 2372
rect 25593 2363 25651 2369
rect 25593 2360 25605 2363
rect 25004 2332 25605 2360
rect 25004 2320 25010 2332
rect 25593 2329 25605 2332
rect 25639 2329 25651 2363
rect 26252 2360 26280 2388
rect 27617 2363 27675 2369
rect 27617 2360 27629 2363
rect 26252 2332 27629 2360
rect 25593 2323 25651 2329
rect 27617 2329 27629 2332
rect 27663 2329 27675 2363
rect 27816 2360 27844 2400
rect 27890 2388 27896 2440
rect 27948 2388 27954 2440
rect 28074 2388 28080 2440
rect 28132 2428 28138 2440
rect 28169 2431 28227 2437
rect 28169 2428 28181 2431
rect 28132 2400 28181 2428
rect 28132 2388 28138 2400
rect 28169 2397 28181 2400
rect 28215 2397 28227 2431
rect 28169 2391 28227 2397
rect 28718 2388 28724 2440
rect 28776 2388 28782 2440
rect 29362 2388 29368 2440
rect 29420 2388 29426 2440
rect 29546 2388 29552 2440
rect 29604 2428 29610 2440
rect 29641 2431 29699 2437
rect 29641 2428 29653 2431
rect 29604 2400 29653 2428
rect 29604 2388 29610 2400
rect 29641 2397 29653 2400
rect 29687 2397 29699 2431
rect 29641 2391 29699 2397
rect 29822 2388 29828 2440
rect 29880 2428 29886 2440
rect 31312 2437 31340 2468
rect 31726 2468 33609 2496
rect 30193 2431 30251 2437
rect 30193 2428 30205 2431
rect 29880 2400 30205 2428
rect 29880 2388 29886 2400
rect 30193 2397 30205 2400
rect 30239 2397 30251 2431
rect 30193 2391 30251 2397
rect 31297 2431 31355 2437
rect 31297 2397 31309 2431
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 30745 2363 30803 2369
rect 30745 2360 30757 2363
rect 27816 2332 30757 2360
rect 27617 2323 27675 2329
rect 30745 2329 30757 2332
rect 30791 2329 30803 2363
rect 30745 2323 30803 2329
rect 31110 2320 31116 2372
rect 31168 2360 31174 2372
rect 31726 2360 31754 2468
rect 33597 2465 33609 2468
rect 33643 2465 33655 2499
rect 33597 2459 33655 2465
rect 34330 2456 34336 2508
rect 34388 2496 34394 2508
rect 34388 2468 36768 2496
rect 34388 2456 34394 2468
rect 31941 2431 31999 2437
rect 31941 2397 31953 2431
rect 31987 2428 31999 2431
rect 31987 2400 32076 2428
rect 31987 2397 31999 2400
rect 31941 2391 31999 2397
rect 31168 2332 31754 2360
rect 32048 2360 32076 2400
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 34517 2431 34575 2437
rect 34517 2428 34529 2431
rect 34204 2400 34529 2428
rect 34204 2388 34210 2400
rect 34517 2397 34529 2400
rect 34563 2397 34575 2431
rect 34517 2391 34575 2397
rect 35897 2431 35955 2437
rect 35897 2397 35909 2431
rect 35943 2428 35955 2431
rect 35986 2428 35992 2440
rect 35943 2400 35992 2428
rect 35943 2397 35955 2400
rect 35897 2391 35955 2397
rect 35986 2388 35992 2400
rect 36044 2388 36050 2440
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36265 2431 36323 2437
rect 36265 2428 36277 2431
rect 36136 2400 36277 2428
rect 36136 2388 36142 2400
rect 36265 2397 36277 2400
rect 36311 2397 36323 2431
rect 36265 2391 36323 2397
rect 36538 2388 36544 2440
rect 36596 2388 36602 2440
rect 36740 2428 36768 2468
rect 36814 2456 36820 2508
rect 36872 2496 36878 2508
rect 36872 2468 37872 2496
rect 36872 2456 36878 2468
rect 36906 2428 36912 2440
rect 36740 2400 36912 2428
rect 36906 2388 36912 2400
rect 36964 2388 36970 2440
rect 36998 2388 37004 2440
rect 37056 2388 37062 2440
rect 37458 2388 37464 2440
rect 37516 2388 37522 2440
rect 37844 2437 37872 2468
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2397 37611 2431
rect 37553 2391 37611 2397
rect 37829 2431 37887 2437
rect 37829 2397 37841 2431
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 38105 2431 38163 2437
rect 38105 2397 38117 2431
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 32122 2360 32128 2372
rect 32048 2332 32128 2360
rect 31168 2320 31174 2332
rect 32122 2320 32128 2332
rect 32180 2320 32186 2372
rect 32214 2320 32220 2372
rect 32272 2320 32278 2372
rect 32398 2320 32404 2372
rect 32456 2360 32462 2372
rect 32769 2363 32827 2369
rect 32769 2360 32781 2363
rect 32456 2332 32781 2360
rect 32456 2320 32462 2332
rect 32769 2329 32781 2332
rect 32815 2329 32827 2363
rect 32769 2323 32827 2329
rect 33318 2320 33324 2372
rect 33376 2320 33382 2372
rect 33870 2320 33876 2372
rect 33928 2320 33934 2372
rect 34790 2320 34796 2372
rect 34848 2320 34854 2372
rect 35342 2320 35348 2372
rect 35400 2320 35406 2372
rect 36446 2320 36452 2372
rect 36504 2360 36510 2372
rect 37568 2360 37596 2391
rect 38120 2360 38148 2391
rect 38378 2388 38384 2440
rect 38436 2388 38442 2440
rect 38654 2388 38660 2440
rect 38712 2388 38718 2440
rect 38948 2437 38976 2536
rect 39117 2533 39129 2567
rect 39163 2533 39175 2567
rect 39117 2527 39175 2533
rect 39853 2567 39911 2573
rect 39853 2533 39865 2567
rect 39899 2564 39911 2567
rect 40512 2564 40540 2592
rect 39899 2536 40540 2564
rect 40681 2567 40739 2573
rect 39899 2533 39911 2536
rect 39853 2527 39911 2533
rect 40681 2533 40693 2567
rect 40727 2533 40739 2567
rect 40681 2527 40739 2533
rect 40957 2567 41015 2573
rect 40957 2533 40969 2567
rect 41003 2564 41015 2567
rect 41003 2536 43024 2564
rect 41003 2533 41015 2536
rect 40957 2527 41015 2533
rect 40696 2496 40724 2527
rect 40696 2468 41460 2496
rect 38933 2431 38991 2437
rect 38933 2397 38945 2431
rect 38979 2397 38991 2431
rect 38933 2391 38991 2397
rect 39114 2388 39120 2440
rect 39172 2428 39178 2440
rect 39393 2431 39451 2437
rect 39393 2428 39405 2431
rect 39172 2400 39405 2428
rect 39172 2388 39178 2400
rect 39393 2397 39405 2400
rect 39439 2397 39451 2431
rect 39393 2391 39451 2397
rect 39666 2388 39672 2440
rect 39724 2388 39730 2440
rect 39758 2388 39764 2440
rect 39816 2428 39822 2440
rect 40037 2431 40095 2437
rect 40037 2428 40049 2431
rect 39816 2400 40049 2428
rect 39816 2388 39822 2400
rect 40037 2397 40049 2400
rect 40083 2397 40095 2431
rect 40037 2391 40095 2397
rect 40310 2388 40316 2440
rect 40368 2388 40374 2440
rect 40402 2388 40408 2440
rect 40460 2428 40466 2440
rect 40589 2431 40647 2437
rect 40589 2428 40601 2431
rect 40460 2400 40601 2428
rect 40460 2388 40466 2400
rect 40589 2397 40601 2400
rect 40635 2397 40647 2431
rect 40589 2391 40647 2397
rect 40862 2388 40868 2440
rect 40920 2388 40926 2440
rect 41432 2437 41460 2468
rect 42996 2437 43024 2536
rect 41141 2431 41199 2437
rect 41141 2397 41153 2431
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 41417 2431 41475 2437
rect 41417 2397 41429 2431
rect 41463 2397 41475 2431
rect 41417 2391 41475 2397
rect 42981 2431 43039 2437
rect 42981 2397 42993 2431
rect 43027 2397 43039 2431
rect 42981 2391 43039 2397
rect 36504 2332 37596 2360
rect 37660 2332 38148 2360
rect 36504 2320 36510 2332
rect 25133 2295 25191 2301
rect 25133 2292 25145 2295
rect 24872 2264 25145 2292
rect 24581 2255 24639 2261
rect 25133 2261 25145 2264
rect 25179 2261 25191 2295
rect 25133 2255 25191 2261
rect 25498 2252 25504 2304
rect 25556 2292 25562 2304
rect 26237 2295 26295 2301
rect 26237 2292 26249 2295
rect 25556 2264 26249 2292
rect 25556 2252 25562 2264
rect 26237 2261 26249 2264
rect 26283 2261 26295 2295
rect 26237 2255 26295 2261
rect 26326 2252 26332 2304
rect 26384 2292 26390 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26384 2264 27169 2292
rect 26384 2252 26390 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 28350 2252 28356 2304
rect 28408 2292 28414 2304
rect 29733 2295 29791 2301
rect 29733 2292 29745 2295
rect 28408 2264 29745 2292
rect 28408 2252 28414 2264
rect 29733 2261 29745 2264
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 30190 2252 30196 2304
rect 30248 2292 30254 2304
rect 31389 2295 31447 2301
rect 31389 2292 31401 2295
rect 30248 2264 31401 2292
rect 30248 2252 30254 2264
rect 31389 2261 31401 2264
rect 31435 2261 31447 2295
rect 31389 2255 31447 2261
rect 31662 2252 31668 2304
rect 31720 2292 31726 2304
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 31720 2264 32321 2292
rect 31720 2252 31726 2264
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 33965 2295 34023 2301
rect 33965 2292 33977 2295
rect 32916 2264 33977 2292
rect 32916 2252 32922 2264
rect 33965 2261 33977 2264
rect 34011 2261 34023 2295
rect 33965 2255 34023 2261
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 34885 2295 34943 2301
rect 34885 2292 34897 2295
rect 34204 2264 34897 2292
rect 34204 2252 34210 2264
rect 34885 2261 34897 2264
rect 34931 2261 34943 2295
rect 34885 2255 34943 2261
rect 34974 2252 34980 2304
rect 35032 2292 35038 2304
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 35032 2264 36369 2292
rect 35032 2252 35038 2264
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 36357 2255 36415 2261
rect 37090 2252 37096 2304
rect 37148 2292 37154 2304
rect 37660 2292 37688 2332
rect 38470 2320 38476 2372
rect 38528 2360 38534 2372
rect 38528 2332 39528 2360
rect 38528 2320 38534 2332
rect 37148 2264 37688 2292
rect 37737 2295 37795 2301
rect 37148 2252 37154 2264
rect 37737 2261 37749 2295
rect 37783 2292 37795 2295
rect 37826 2292 37832 2304
rect 37783 2264 37832 2292
rect 37783 2261 37795 2264
rect 37737 2255 37795 2261
rect 37826 2252 37832 2264
rect 37884 2252 37890 2304
rect 38010 2252 38016 2304
rect 38068 2252 38074 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38562 2252 38568 2304
rect 38620 2252 38626 2304
rect 38841 2295 38899 2301
rect 38841 2261 38853 2295
rect 38887 2292 38899 2295
rect 38930 2292 38936 2304
rect 38887 2264 38936 2292
rect 38887 2261 38899 2264
rect 38841 2255 38899 2261
rect 38930 2252 38936 2264
rect 38988 2252 38994 2304
rect 39500 2301 39528 2332
rect 39942 2320 39948 2372
rect 40000 2360 40006 2372
rect 41156 2360 41184 2391
rect 40000 2332 41184 2360
rect 40000 2320 40006 2332
rect 39485 2295 39543 2301
rect 39485 2261 39497 2295
rect 39531 2261 39543 2295
rect 39485 2255 39543 2261
rect 1104 2202 44040 2224
rect 1104 2150 11644 2202
rect 11696 2150 11708 2202
rect 11760 2150 11772 2202
rect 11824 2150 11836 2202
rect 11888 2150 11900 2202
rect 11952 2150 22338 2202
rect 22390 2150 22402 2202
rect 22454 2150 22466 2202
rect 22518 2150 22530 2202
rect 22582 2150 22594 2202
rect 22646 2150 33032 2202
rect 33084 2150 33096 2202
rect 33148 2150 33160 2202
rect 33212 2150 33224 2202
rect 33276 2150 33288 2202
rect 33340 2150 43726 2202
rect 43778 2150 43790 2202
rect 43842 2150 43854 2202
rect 43906 2150 43918 2202
rect 43970 2150 43982 2202
rect 44034 2150 44040 2202
rect 1104 2128 44040 2150
rect 4890 2048 4896 2100
rect 4948 2048 4954 2100
rect 5534 2048 5540 2100
rect 5592 2048 5598 2100
rect 5902 2048 5908 2100
rect 5960 2088 5966 2100
rect 10870 2088 10876 2100
rect 5960 2060 10876 2088
rect 5960 2048 5966 2060
rect 10870 2048 10876 2060
rect 10928 2048 10934 2100
rect 11422 2048 11428 2100
rect 11480 2088 11486 2100
rect 19426 2088 19432 2100
rect 11480 2060 19432 2088
rect 11480 2048 11486 2060
rect 19426 2048 19432 2060
rect 19484 2048 19490 2100
rect 20806 2048 20812 2100
rect 20864 2048 20870 2100
rect 20990 2048 20996 2100
rect 21048 2088 21054 2100
rect 32398 2088 32404 2100
rect 21048 2060 32404 2088
rect 21048 2048 21054 2060
rect 32398 2048 32404 2060
rect 32456 2048 32462 2100
rect 38286 2088 38292 2100
rect 35866 2060 38292 2088
rect 4908 1748 4936 2048
rect 5552 2020 5580 2048
rect 11054 2020 11060 2032
rect 5552 1992 11060 2020
rect 11054 1980 11060 1992
rect 11112 1980 11118 2032
rect 15194 2020 15200 2032
rect 11256 1992 15200 2020
rect 7926 1912 7932 1964
rect 7984 1912 7990 1964
rect 8294 1912 8300 1964
rect 8352 1952 8358 1964
rect 11256 1952 11284 1992
rect 15194 1980 15200 1992
rect 15252 1980 15258 2032
rect 16942 1980 16948 2032
rect 17000 2020 17006 2032
rect 20824 2020 20852 2048
rect 26786 2020 26792 2032
rect 17000 1992 20852 2020
rect 20916 1992 26792 2020
rect 17000 1980 17006 1992
rect 8352 1924 11284 1952
rect 8352 1912 8358 1924
rect 11330 1912 11336 1964
rect 11388 1952 11394 1964
rect 11388 1924 18000 1952
rect 11388 1912 11394 1924
rect 7944 1884 7972 1912
rect 13814 1884 13820 1896
rect 7944 1856 13820 1884
rect 13814 1844 13820 1856
rect 13872 1844 13878 1896
rect 17678 1844 17684 1896
rect 17736 1844 17742 1896
rect 17696 1816 17724 1844
rect 12360 1788 17724 1816
rect 17972 1816 18000 1924
rect 18046 1844 18052 1896
rect 18104 1884 18110 1896
rect 20916 1884 20944 1992
rect 26786 1980 26792 1992
rect 26844 1980 26850 2032
rect 29362 1980 29368 2032
rect 29420 1980 29426 2032
rect 30374 1980 30380 2032
rect 30432 2020 30438 2032
rect 32214 2020 32220 2032
rect 30432 1992 32220 2020
rect 30432 1980 30438 1992
rect 32214 1980 32220 1992
rect 32272 1980 32278 2032
rect 29380 1952 29408 1980
rect 35866 1952 35894 2060
rect 38286 2048 38292 2060
rect 38344 2048 38350 2100
rect 38470 2048 38476 2100
rect 38528 2048 38534 2100
rect 38562 2048 38568 2100
rect 38620 2048 38626 2100
rect 18104 1856 20944 1884
rect 21008 1924 29408 1952
rect 31726 1924 35894 1952
rect 18104 1844 18110 1856
rect 21008 1816 21036 1924
rect 21542 1844 21548 1896
rect 21600 1844 21606 1896
rect 31726 1884 31754 1924
rect 22066 1856 31754 1884
rect 17972 1788 21036 1816
rect 12158 1748 12164 1760
rect 4908 1720 12164 1748
rect 12158 1708 12164 1720
rect 12216 1708 12222 1760
rect 6546 1640 6552 1692
rect 6604 1640 6610 1692
rect 7374 1640 7380 1692
rect 7432 1640 7438 1692
rect 8202 1640 8208 1692
rect 8260 1680 8266 1692
rect 12360 1680 12388 1788
rect 21560 1748 21588 1844
rect 21910 1776 21916 1828
rect 21968 1816 21974 1828
rect 22066 1816 22094 1856
rect 32122 1844 32128 1896
rect 32180 1884 32186 1896
rect 38488 1884 38516 2048
rect 32180 1856 38516 1884
rect 32180 1844 32186 1856
rect 21968 1788 22094 1816
rect 21968 1776 21974 1788
rect 23014 1776 23020 1828
rect 23072 1816 23078 1828
rect 38580 1816 38608 2048
rect 23072 1788 38608 1816
rect 23072 1776 23078 1788
rect 8260 1652 12388 1680
rect 12452 1720 21588 1748
rect 8260 1640 8266 1652
rect 6564 1476 6592 1640
rect 7392 1612 7420 1640
rect 12452 1612 12480 1720
rect 31386 1708 31392 1760
rect 31444 1748 31450 1760
rect 34974 1748 34980 1760
rect 31444 1720 34980 1748
rect 31444 1708 31450 1720
rect 34974 1708 34980 1720
rect 35032 1708 35038 1760
rect 35066 1708 35072 1760
rect 35124 1748 35130 1760
rect 36998 1748 37004 1760
rect 35124 1720 37004 1748
rect 35124 1708 35130 1720
rect 36998 1708 37004 1720
rect 37056 1708 37062 1760
rect 12802 1640 12808 1692
rect 12860 1680 12866 1692
rect 26418 1680 26424 1692
rect 12860 1652 26424 1680
rect 12860 1640 12866 1652
rect 26418 1640 26424 1652
rect 26476 1640 26482 1692
rect 7392 1584 12480 1612
rect 16666 1572 16672 1624
rect 16724 1612 16730 1624
rect 19150 1612 19156 1624
rect 16724 1584 19156 1612
rect 16724 1572 16730 1584
rect 19150 1572 19156 1584
rect 19208 1572 19214 1624
rect 38286 1572 38292 1624
rect 38344 1612 38350 1624
rect 39666 1612 39672 1624
rect 38344 1584 39672 1612
rect 38344 1572 38350 1584
rect 39666 1572 39672 1584
rect 39724 1572 39730 1624
rect 8570 1504 8576 1556
rect 8628 1544 8634 1556
rect 9306 1544 9312 1556
rect 8628 1516 9312 1544
rect 8628 1504 8634 1516
rect 9306 1504 9312 1516
rect 9364 1504 9370 1556
rect 17126 1504 17132 1556
rect 17184 1544 17190 1556
rect 23198 1544 23204 1556
rect 17184 1516 23204 1544
rect 17184 1504 17190 1516
rect 23198 1504 23204 1516
rect 23256 1504 23262 1556
rect 34422 1504 34428 1556
rect 34480 1544 34486 1556
rect 36538 1544 36544 1556
rect 34480 1516 36544 1544
rect 34480 1504 34486 1516
rect 36538 1504 36544 1516
rect 36596 1504 36602 1556
rect 37458 1504 37464 1556
rect 37516 1504 37522 1556
rect 38470 1504 38476 1556
rect 38528 1544 38534 1556
rect 39758 1544 39764 1556
rect 38528 1516 39764 1544
rect 38528 1504 38534 1516
rect 39758 1504 39764 1516
rect 39816 1504 39822 1556
rect 23750 1476 23756 1488
rect 6564 1448 23756 1476
rect 23750 1436 23756 1448
rect 23808 1436 23814 1488
rect 31846 1436 31852 1488
rect 31904 1476 31910 1488
rect 32858 1476 32864 1488
rect 31904 1448 32864 1476
rect 31904 1436 31910 1448
rect 32858 1436 32864 1448
rect 32916 1436 32922 1488
rect 35618 1436 35624 1488
rect 35676 1476 35682 1488
rect 37476 1476 37504 1504
rect 35676 1448 37504 1476
rect 35676 1436 35682 1448
rect 38562 1436 38568 1488
rect 38620 1476 38626 1488
rect 40310 1476 40316 1488
rect 38620 1448 40316 1476
rect 38620 1436 38626 1448
rect 40310 1436 40316 1448
rect 40368 1436 40374 1488
rect 5626 1368 5632 1420
rect 5684 1408 5690 1420
rect 6270 1408 6276 1420
rect 5684 1380 6276 1408
rect 5684 1368 5690 1380
rect 6270 1368 6276 1380
rect 6328 1368 6334 1420
rect 6822 1368 6828 1420
rect 6880 1408 6886 1420
rect 6880 1380 9628 1408
rect 6880 1368 6886 1380
rect 9600 1068 9628 1380
rect 11146 1368 11152 1420
rect 11204 1408 11210 1420
rect 11790 1408 11796 1420
rect 11204 1380 11796 1408
rect 11204 1368 11210 1380
rect 11790 1368 11796 1380
rect 11848 1368 11854 1420
rect 12710 1368 12716 1420
rect 12768 1408 12774 1420
rect 13170 1408 13176 1420
rect 12768 1380 13176 1408
rect 12768 1368 12774 1380
rect 13170 1368 13176 1380
rect 13228 1368 13234 1420
rect 32398 1368 32404 1420
rect 32456 1408 32462 1420
rect 34146 1408 34152 1420
rect 32456 1380 34152 1408
rect 32456 1368 32462 1380
rect 34146 1368 34152 1380
rect 34204 1368 34210 1420
rect 37090 1368 37096 1420
rect 37148 1408 37154 1420
rect 38378 1408 38384 1420
rect 37148 1380 38384 1408
rect 37148 1368 37154 1380
rect 38378 1368 38384 1380
rect 38436 1368 38442 1420
rect 39666 1368 39672 1420
rect 39724 1408 39730 1420
rect 40862 1408 40868 1420
rect 39724 1380 40868 1408
rect 39724 1368 39730 1380
rect 40862 1368 40868 1380
rect 40920 1368 40926 1420
rect 15102 1300 15108 1352
rect 15160 1340 15166 1352
rect 35342 1340 35348 1352
rect 15160 1312 35348 1340
rect 15160 1300 15166 1312
rect 35342 1300 35348 1312
rect 35400 1300 35406 1352
rect 15562 1232 15568 1284
rect 15620 1272 15626 1284
rect 33778 1272 33784 1284
rect 15620 1244 33784 1272
rect 15620 1232 15626 1244
rect 33778 1232 33784 1244
rect 33836 1232 33842 1284
rect 16114 1164 16120 1216
rect 16172 1204 16178 1216
rect 33686 1204 33692 1216
rect 16172 1176 33692 1204
rect 16172 1164 16178 1176
rect 33686 1164 33692 1176
rect 33744 1164 33750 1216
rect 15838 1096 15844 1148
rect 15896 1136 15902 1148
rect 32030 1136 32036 1148
rect 15896 1108 32036 1136
rect 15896 1096 15902 1108
rect 32030 1096 32036 1108
rect 32088 1096 32094 1148
rect 9600 1040 16574 1068
rect 16546 1000 16574 1040
rect 17494 1028 17500 1080
rect 17552 1068 17558 1080
rect 33870 1068 33876 1080
rect 17552 1040 33876 1068
rect 17552 1028 17558 1040
rect 33870 1028 33876 1040
rect 33928 1028 33934 1080
rect 23842 1000 23848 1012
rect 16546 972 23848 1000
rect 23842 960 23848 972
rect 23900 960 23906 1012
rect 10870 892 10876 944
rect 10928 932 10934 944
rect 20070 932 20076 944
rect 10928 904 20076 932
rect 10928 892 10934 904
rect 20070 892 20076 904
rect 20128 892 20134 944
<< via1 >>
rect 22192 7760 22244 7812
rect 31392 7760 31444 7812
rect 19064 7692 19116 7744
rect 35900 7692 35952 7744
rect 11644 7590 11696 7642
rect 11708 7590 11760 7642
rect 11772 7590 11824 7642
rect 11836 7590 11888 7642
rect 11900 7590 11952 7642
rect 22338 7590 22390 7642
rect 22402 7590 22454 7642
rect 22466 7590 22518 7642
rect 22530 7590 22582 7642
rect 22594 7590 22646 7642
rect 33032 7590 33084 7642
rect 33096 7590 33148 7642
rect 33160 7590 33212 7642
rect 33224 7590 33276 7642
rect 33288 7590 33340 7642
rect 43726 7590 43778 7642
rect 43790 7590 43842 7642
rect 43854 7590 43906 7642
rect 43918 7590 43970 7642
rect 43982 7590 44034 7642
rect 1308 7488 1360 7540
rect 3792 7488 3844 7540
rect 5540 7488 5592 7540
rect 7656 7488 7708 7540
rect 9772 7488 9824 7540
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 14004 7488 14056 7540
rect 16580 7488 16632 7540
rect 4068 7352 4120 7404
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 16764 7395 16816 7404
rect 16764 7361 16773 7395
rect 16773 7361 16807 7395
rect 16807 7361 16816 7395
rect 16764 7352 16816 7361
rect 21088 7488 21140 7540
rect 20720 7420 20772 7472
rect 22836 7488 22888 7540
rect 24676 7488 24728 7540
rect 26700 7488 26752 7540
rect 28908 7488 28960 7540
rect 30932 7488 30984 7540
rect 32956 7488 33008 7540
rect 35164 7488 35216 7540
rect 37280 7488 37332 7540
rect 18604 7352 18656 7404
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 21916 7352 21968 7404
rect 23388 7352 23440 7404
rect 23480 7395 23532 7404
rect 23480 7361 23489 7395
rect 23489 7361 23523 7395
rect 23523 7361 23532 7395
rect 23480 7352 23532 7361
rect 24860 7352 24912 7404
rect 26884 7352 26936 7404
rect 29000 7395 29052 7404
rect 29000 7361 29009 7395
rect 29009 7361 29043 7395
rect 29043 7361 29052 7395
rect 29000 7352 29052 7361
rect 31760 7352 31812 7404
rect 39672 7488 39724 7540
rect 41512 7488 41564 7540
rect 43628 7488 43680 7540
rect 34336 7284 34388 7336
rect 35348 7395 35400 7404
rect 35348 7361 35357 7395
rect 35357 7361 35391 7395
rect 35391 7361 35400 7395
rect 35348 7352 35400 7361
rect 35532 7284 35584 7336
rect 22192 7216 22244 7268
rect 17316 7148 17368 7200
rect 18236 7148 18288 7200
rect 18604 7148 18656 7200
rect 40224 7352 40276 7404
rect 41696 7395 41748 7404
rect 41696 7361 41705 7395
rect 41705 7361 41739 7395
rect 41739 7361 41748 7395
rect 41696 7352 41748 7361
rect 43168 7395 43220 7404
rect 43168 7361 43177 7395
rect 43177 7361 43211 7395
rect 43211 7361 43220 7395
rect 43168 7352 43220 7361
rect 40500 7284 40552 7336
rect 40040 7216 40092 7268
rect 6297 7046 6349 7098
rect 6361 7046 6413 7098
rect 6425 7046 6477 7098
rect 6489 7046 6541 7098
rect 6553 7046 6605 7098
rect 16991 7046 17043 7098
rect 17055 7046 17107 7098
rect 17119 7046 17171 7098
rect 17183 7046 17235 7098
rect 17247 7046 17299 7098
rect 27685 7046 27737 7098
rect 27749 7046 27801 7098
rect 27813 7046 27865 7098
rect 27877 7046 27929 7098
rect 27941 7046 27993 7098
rect 38379 7046 38431 7098
rect 38443 7046 38495 7098
rect 38507 7046 38559 7098
rect 38571 7046 38623 7098
rect 38635 7046 38687 7098
rect 17316 6944 17368 6996
rect 21088 6944 21140 6996
rect 23388 6944 23440 6996
rect 36728 6944 36780 6996
rect 26884 6876 26936 6928
rect 34428 6876 34480 6928
rect 23020 6783 23072 6792
rect 23020 6749 23029 6783
rect 23029 6749 23063 6783
rect 23063 6749 23072 6783
rect 23020 6740 23072 6749
rect 23480 6740 23532 6792
rect 11644 6502 11696 6554
rect 11708 6502 11760 6554
rect 11772 6502 11824 6554
rect 11836 6502 11888 6554
rect 11900 6502 11952 6554
rect 22338 6502 22390 6554
rect 22402 6502 22454 6554
rect 22466 6502 22518 6554
rect 22530 6502 22582 6554
rect 22594 6502 22646 6554
rect 33032 6502 33084 6554
rect 33096 6502 33148 6554
rect 33160 6502 33212 6554
rect 33224 6502 33276 6554
rect 33288 6502 33340 6554
rect 43726 6502 43778 6554
rect 43790 6502 43842 6554
rect 43854 6502 43906 6554
rect 43918 6502 43970 6554
rect 43982 6502 44034 6554
rect 5724 6196 5776 6248
rect 35808 6196 35860 6248
rect 4068 6128 4120 6180
rect 33600 6128 33652 6180
rect 6297 5958 6349 6010
rect 6361 5958 6413 6010
rect 6425 5958 6477 6010
rect 6489 5958 6541 6010
rect 6553 5958 6605 6010
rect 16991 5958 17043 6010
rect 17055 5958 17107 6010
rect 17119 5958 17171 6010
rect 17183 5958 17235 6010
rect 17247 5958 17299 6010
rect 27685 5958 27737 6010
rect 27749 5958 27801 6010
rect 27813 5958 27865 6010
rect 27877 5958 27929 6010
rect 27941 5958 27993 6010
rect 38379 5958 38431 6010
rect 38443 5958 38495 6010
rect 38507 5958 38559 6010
rect 38571 5958 38623 6010
rect 38635 5958 38687 6010
rect 16764 5856 16816 5908
rect 24860 5899 24912 5908
rect 24860 5865 24869 5899
rect 24869 5865 24903 5899
rect 24903 5865 24912 5899
rect 24860 5856 24912 5865
rect 16488 5652 16540 5704
rect 38936 5652 38988 5704
rect 35900 5516 35952 5568
rect 38016 5516 38068 5568
rect 11644 5414 11696 5466
rect 11708 5414 11760 5466
rect 11772 5414 11824 5466
rect 11836 5414 11888 5466
rect 11900 5414 11952 5466
rect 22338 5414 22390 5466
rect 22402 5414 22454 5466
rect 22466 5414 22518 5466
rect 22530 5414 22582 5466
rect 22594 5414 22646 5466
rect 33032 5414 33084 5466
rect 33096 5414 33148 5466
rect 33160 5414 33212 5466
rect 33224 5414 33276 5466
rect 33288 5414 33340 5466
rect 43726 5414 43778 5466
rect 43790 5414 43842 5466
rect 43854 5414 43906 5466
rect 43918 5414 43970 5466
rect 43982 5414 44034 5466
rect 6297 4870 6349 4922
rect 6361 4870 6413 4922
rect 6425 4870 6477 4922
rect 6489 4870 6541 4922
rect 6553 4870 6605 4922
rect 16991 4870 17043 4922
rect 17055 4870 17107 4922
rect 17119 4870 17171 4922
rect 17183 4870 17235 4922
rect 17247 4870 17299 4922
rect 27685 4870 27737 4922
rect 27749 4870 27801 4922
rect 27813 4870 27865 4922
rect 27877 4870 27929 4922
rect 27941 4870 27993 4922
rect 38379 4870 38431 4922
rect 38443 4870 38495 4922
rect 38507 4870 38559 4922
rect 38571 4870 38623 4922
rect 38635 4870 38687 4922
rect 9680 4700 9732 4752
rect 19432 4700 19484 4752
rect 10232 4632 10284 4684
rect 28816 4632 28868 4684
rect 6184 4564 6236 4616
rect 24216 4564 24268 4616
rect 14096 4496 14148 4548
rect 25964 4496 26016 4548
rect 8668 4428 8720 4480
rect 24492 4428 24544 4480
rect 11644 4326 11696 4378
rect 11708 4326 11760 4378
rect 11772 4326 11824 4378
rect 11836 4326 11888 4378
rect 11900 4326 11952 4378
rect 22338 4326 22390 4378
rect 22402 4326 22454 4378
rect 22466 4326 22518 4378
rect 22530 4326 22582 4378
rect 22594 4326 22646 4378
rect 33032 4326 33084 4378
rect 33096 4326 33148 4378
rect 33160 4326 33212 4378
rect 33224 4326 33276 4378
rect 33288 4326 33340 4378
rect 43726 4326 43778 4378
rect 43790 4326 43842 4378
rect 43854 4326 43906 4378
rect 43918 4326 43970 4378
rect 43982 4326 44034 4378
rect 14464 4224 14516 4276
rect 25504 4224 25556 4276
rect 13912 4156 13964 4208
rect 33416 4156 33468 4208
rect 13912 4020 13964 4072
rect 10324 3952 10376 4004
rect 9956 3884 10008 3936
rect 20168 3884 20220 3936
rect 21732 3884 21784 3936
rect 25412 3884 25464 3936
rect 26240 3884 26292 3936
rect 30012 3884 30064 3936
rect 6297 3782 6349 3834
rect 6361 3782 6413 3834
rect 6425 3782 6477 3834
rect 6489 3782 6541 3834
rect 6553 3782 6605 3834
rect 16991 3782 17043 3834
rect 17055 3782 17107 3834
rect 17119 3782 17171 3834
rect 17183 3782 17235 3834
rect 17247 3782 17299 3834
rect 27685 3782 27737 3834
rect 27749 3782 27801 3834
rect 27813 3782 27865 3834
rect 27877 3782 27929 3834
rect 27941 3782 27993 3834
rect 38379 3782 38431 3834
rect 38443 3782 38495 3834
rect 38507 3782 38559 3834
rect 38571 3782 38623 3834
rect 38635 3782 38687 3834
rect 15108 3680 15160 3732
rect 16672 3612 16724 3664
rect 23480 3612 23532 3664
rect 9312 3544 9364 3596
rect 16764 3476 16816 3528
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 18420 3476 18472 3528
rect 18604 3408 18656 3460
rect 19248 3476 19300 3528
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 19432 3408 19484 3460
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 22100 3544 22152 3596
rect 21732 3476 21784 3528
rect 22008 3476 22060 3528
rect 23204 3519 23256 3528
rect 23204 3485 23213 3519
rect 23213 3485 23247 3519
rect 23247 3485 23256 3519
rect 23204 3476 23256 3485
rect 23848 3476 23900 3528
rect 27068 3680 27120 3732
rect 25688 3612 25740 3664
rect 27988 3612 28040 3664
rect 24952 3544 25004 3596
rect 29000 3680 29052 3732
rect 33600 3723 33652 3732
rect 33600 3689 33609 3723
rect 33609 3689 33643 3723
rect 33643 3689 33652 3723
rect 33600 3680 33652 3689
rect 29828 3612 29880 3664
rect 16304 3340 16356 3392
rect 17776 3340 17828 3392
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 19340 3383 19392 3392
rect 19340 3349 19349 3383
rect 19349 3349 19383 3383
rect 19383 3349 19392 3383
rect 19340 3340 19392 3349
rect 19708 3383 19760 3392
rect 19708 3349 19717 3383
rect 19717 3349 19751 3383
rect 19751 3349 19760 3383
rect 19708 3340 19760 3349
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 20812 3340 20864 3392
rect 20904 3383 20956 3392
rect 20904 3349 20913 3383
rect 20913 3349 20947 3383
rect 20947 3349 20956 3383
rect 20904 3340 20956 3349
rect 21180 3383 21232 3392
rect 21180 3349 21189 3383
rect 21189 3349 21223 3383
rect 21223 3349 21232 3383
rect 21180 3340 21232 3349
rect 21456 3383 21508 3392
rect 21456 3349 21465 3383
rect 21465 3349 21499 3383
rect 21499 3349 21508 3383
rect 21456 3340 21508 3349
rect 23664 3408 23716 3460
rect 25412 3519 25464 3528
rect 25412 3485 25421 3519
rect 25421 3485 25455 3519
rect 25455 3485 25464 3519
rect 25412 3476 25464 3485
rect 25504 3476 25556 3528
rect 25964 3519 26016 3528
rect 25964 3485 25973 3519
rect 25973 3485 26007 3519
rect 26007 3485 26016 3519
rect 25964 3476 26016 3485
rect 26240 3519 26292 3528
rect 26240 3485 26249 3519
rect 26249 3485 26283 3519
rect 26283 3485 26292 3519
rect 26240 3476 26292 3485
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 26792 3519 26844 3528
rect 26792 3485 26801 3519
rect 26801 3485 26835 3519
rect 26835 3485 26844 3519
rect 26792 3476 26844 3485
rect 29552 3544 29604 3596
rect 27160 3476 27212 3528
rect 27620 3476 27672 3528
rect 28264 3519 28316 3528
rect 28264 3485 28273 3519
rect 28273 3485 28307 3519
rect 28307 3485 28316 3519
rect 28264 3476 28316 3485
rect 28540 3519 28592 3528
rect 28540 3485 28549 3519
rect 28549 3485 28583 3519
rect 28583 3485 28592 3519
rect 28540 3476 28592 3485
rect 28816 3519 28868 3528
rect 28816 3485 28825 3519
rect 28825 3485 28859 3519
rect 28859 3485 28868 3519
rect 28816 3476 28868 3485
rect 36820 3476 36872 3528
rect 22008 3383 22060 3392
rect 22008 3349 22017 3383
rect 22017 3349 22051 3383
rect 22051 3349 22060 3383
rect 22008 3340 22060 3349
rect 22192 3340 22244 3392
rect 22928 3340 22980 3392
rect 23940 3340 23992 3392
rect 24400 3383 24452 3392
rect 24400 3349 24409 3383
rect 24409 3349 24443 3383
rect 24443 3349 24452 3383
rect 24400 3340 24452 3349
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 26700 3408 26752 3460
rect 26148 3340 26200 3392
rect 26332 3383 26384 3392
rect 26332 3349 26341 3383
rect 26341 3349 26375 3383
rect 26375 3349 26384 3383
rect 26332 3340 26384 3349
rect 26884 3383 26936 3392
rect 26884 3349 26893 3383
rect 26893 3349 26927 3383
rect 26927 3349 26936 3383
rect 26884 3340 26936 3349
rect 28724 3408 28776 3460
rect 32036 3408 32088 3460
rect 33508 3451 33560 3460
rect 33508 3417 33517 3451
rect 33517 3417 33551 3451
rect 33551 3417 33560 3451
rect 33508 3408 33560 3417
rect 28080 3383 28132 3392
rect 28080 3349 28089 3383
rect 28089 3349 28123 3383
rect 28123 3349 28132 3383
rect 28080 3340 28132 3349
rect 28632 3383 28684 3392
rect 28632 3349 28641 3383
rect 28641 3349 28675 3383
rect 28675 3349 28684 3383
rect 28632 3340 28684 3349
rect 32772 3340 32824 3392
rect 34980 3340 35032 3392
rect 36912 3340 36964 3392
rect 11644 3238 11696 3290
rect 11708 3238 11760 3290
rect 11772 3238 11824 3290
rect 11836 3238 11888 3290
rect 11900 3238 11952 3290
rect 22338 3238 22390 3290
rect 22402 3238 22454 3290
rect 22466 3238 22518 3290
rect 22530 3238 22582 3290
rect 22594 3238 22646 3290
rect 33032 3238 33084 3290
rect 33096 3238 33148 3290
rect 33160 3238 33212 3290
rect 33224 3238 33276 3290
rect 33288 3238 33340 3290
rect 43726 3238 43778 3290
rect 43790 3238 43842 3290
rect 43854 3238 43906 3290
rect 43918 3238 43970 3290
rect 43982 3238 44034 3290
rect 9312 3179 9364 3188
rect 9312 3145 9321 3179
rect 9321 3145 9355 3179
rect 9355 3145 9364 3179
rect 9312 3136 9364 3145
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 18052 3068 18104 3120
rect 19156 3179 19208 3188
rect 19156 3145 19165 3179
rect 19165 3145 19199 3179
rect 19199 3145 19208 3179
rect 19156 3136 19208 3145
rect 19340 3136 19392 3188
rect 19984 3136 20036 3188
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 14004 3000 14056 3052
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14648 3043 14700 3052
rect 14648 3009 14657 3043
rect 14657 3009 14691 3043
rect 14691 3009 14700 3043
rect 14648 3000 14700 3009
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 16212 3043 16264 3052
rect 16212 3009 16221 3043
rect 16221 3009 16255 3043
rect 16255 3009 16264 3043
rect 16212 3000 16264 3009
rect 16488 3043 16540 3052
rect 16488 3009 16497 3043
rect 16497 3009 16531 3043
rect 16531 3009 16540 3043
rect 16488 3000 16540 3009
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 13820 2932 13872 2984
rect 14096 2932 14148 2984
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 15016 2864 15068 2916
rect 15108 2839 15160 2848
rect 15108 2805 15117 2839
rect 15117 2805 15151 2839
rect 15151 2805 15160 2839
rect 15108 2796 15160 2805
rect 15292 2796 15344 2848
rect 15568 2796 15620 2848
rect 15844 2796 15896 2848
rect 16120 2796 16172 2848
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 18788 3000 18840 3052
rect 20812 3136 20864 3188
rect 21456 3136 21508 3188
rect 22008 3136 22060 3188
rect 22928 3136 22980 3188
rect 24400 3068 24452 3120
rect 25228 3136 25280 3188
rect 26332 3136 26384 3188
rect 19616 3043 19668 3052
rect 19616 3009 19625 3043
rect 19625 3009 19659 3043
rect 19659 3009 19668 3043
rect 19616 3000 19668 3009
rect 19892 3000 19944 3052
rect 20812 3000 20864 3052
rect 23756 3000 23808 3052
rect 24216 3043 24268 3052
rect 24216 3009 24225 3043
rect 24225 3009 24259 3043
rect 24259 3009 24268 3043
rect 24216 3000 24268 3009
rect 24492 3043 24544 3052
rect 24492 3009 24501 3043
rect 24501 3009 24535 3043
rect 24535 3009 24544 3043
rect 24492 3000 24544 3009
rect 26240 3000 26292 3052
rect 26700 3068 26752 3120
rect 26884 3068 26936 3120
rect 28080 3136 28132 3188
rect 28632 3136 28684 3188
rect 30564 3136 30616 3188
rect 33048 3136 33100 3188
rect 34520 3136 34572 3188
rect 35532 3136 35584 3188
rect 35624 3136 35676 3188
rect 28908 3000 28960 3052
rect 29000 3000 29052 3052
rect 33416 3068 33468 3120
rect 34980 3111 35032 3120
rect 34980 3077 34989 3111
rect 34989 3077 35023 3111
rect 35023 3077 35032 3111
rect 34980 3068 35032 3077
rect 35256 3068 35308 3120
rect 30012 3000 30064 3052
rect 18328 2907 18380 2916
rect 18328 2873 18337 2907
rect 18337 2873 18371 2907
rect 18371 2873 18380 2907
rect 18328 2864 18380 2873
rect 19340 2932 19392 2984
rect 23572 2932 23624 2984
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 17500 2796 17552 2848
rect 18880 2839 18932 2848
rect 18880 2805 18889 2839
rect 18889 2805 18923 2839
rect 18923 2805 18932 2839
rect 18880 2796 18932 2805
rect 19800 2907 19852 2916
rect 19800 2873 19809 2907
rect 19809 2873 19843 2907
rect 19843 2873 19852 2907
rect 19800 2864 19852 2873
rect 20996 2864 21048 2916
rect 22008 2864 22060 2916
rect 20260 2839 20312 2848
rect 20260 2805 20269 2839
rect 20269 2805 20303 2839
rect 20303 2805 20312 2839
rect 20260 2796 20312 2805
rect 20628 2796 20680 2848
rect 21364 2839 21416 2848
rect 21364 2805 21373 2839
rect 21373 2805 21407 2839
rect 21407 2805 21416 2839
rect 21364 2796 21416 2805
rect 22100 2796 22152 2848
rect 22836 2839 22888 2848
rect 22836 2805 22845 2839
rect 22845 2805 22879 2839
rect 22879 2805 22888 2839
rect 22836 2796 22888 2805
rect 23112 2796 23164 2848
rect 24860 2932 24912 2984
rect 29092 2932 29144 2984
rect 32312 3000 32364 3052
rect 33692 3000 33744 3052
rect 33784 3000 33836 3052
rect 35348 3043 35400 3052
rect 35348 3009 35357 3043
rect 35357 3009 35391 3043
rect 35391 3009 35400 3043
rect 35348 3000 35400 3009
rect 36820 3068 36872 3120
rect 34704 2932 34756 2984
rect 35716 2932 35768 2984
rect 24952 2864 25004 2916
rect 26976 2864 27028 2916
rect 24492 2796 24544 2848
rect 25044 2796 25096 2848
rect 25596 2796 25648 2848
rect 26056 2796 26108 2848
rect 26608 2796 26660 2848
rect 27528 2864 27580 2916
rect 29736 2864 29788 2916
rect 28356 2796 28408 2848
rect 28908 2796 28960 2848
rect 29460 2796 29512 2848
rect 30288 2864 30340 2916
rect 31944 2864 31996 2916
rect 32312 2839 32364 2848
rect 32312 2805 32321 2839
rect 32321 2805 32355 2839
rect 32355 2805 32364 2839
rect 32312 2796 32364 2805
rect 32496 2864 32548 2916
rect 33600 2864 33652 2916
rect 35992 2864 36044 2916
rect 37740 3000 37792 3052
rect 38844 3000 38896 3052
rect 39396 3043 39448 3052
rect 39396 3009 39405 3043
rect 39405 3009 39439 3043
rect 39439 3009 39448 3043
rect 39396 3000 39448 3009
rect 40132 2932 40184 2984
rect 36084 2796 36136 2848
rect 36360 2839 36412 2848
rect 36360 2805 36369 2839
rect 36369 2805 36403 2839
rect 36403 2805 36412 2839
rect 36360 2796 36412 2805
rect 37188 2796 37240 2848
rect 38752 2796 38804 2848
rect 39120 2796 39172 2848
rect 40408 2796 40460 2848
rect 6297 2694 6349 2746
rect 6361 2694 6413 2746
rect 6425 2694 6477 2746
rect 6489 2694 6541 2746
rect 6553 2694 6605 2746
rect 16991 2694 17043 2746
rect 17055 2694 17107 2746
rect 17119 2694 17171 2746
rect 17183 2694 17235 2746
rect 17247 2694 17299 2746
rect 27685 2694 27737 2746
rect 27749 2694 27801 2746
rect 27813 2694 27865 2746
rect 27877 2694 27929 2746
rect 27941 2694 27993 2746
rect 38379 2694 38431 2746
rect 38443 2694 38495 2746
rect 38507 2694 38559 2746
rect 38571 2694 38623 2746
rect 38635 2694 38687 2746
rect 5908 2524 5960 2576
rect 6184 2567 6236 2576
rect 6184 2533 6193 2567
rect 6193 2533 6227 2567
rect 6227 2533 6236 2567
rect 6184 2524 6236 2533
rect 6552 2592 6604 2644
rect 8668 2592 8720 2644
rect 5540 2456 5592 2508
rect 4988 2320 5040 2372
rect 5816 2456 5868 2508
rect 6276 2456 6328 2508
rect 6736 2456 6788 2508
rect 8300 2524 8352 2576
rect 9220 2592 9272 2644
rect 9404 2635 9456 2644
rect 9404 2601 9413 2635
rect 9413 2601 9447 2635
rect 9447 2601 9456 2635
rect 9404 2592 9456 2601
rect 9956 2635 10008 2644
rect 9956 2601 9965 2635
rect 9965 2601 9999 2635
rect 9999 2601 10008 2635
rect 9956 2592 10008 2601
rect 10232 2635 10284 2644
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 13268 2592 13320 2644
rect 8760 2456 8812 2508
rect 5264 2320 5316 2372
rect 4896 2252 4948 2304
rect 5540 2252 5592 2304
rect 5632 2252 5684 2304
rect 6552 2388 6604 2440
rect 7012 2320 7064 2372
rect 7380 2388 7432 2440
rect 7656 2388 7708 2440
rect 7932 2388 7984 2440
rect 7288 2320 7340 2372
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 6828 2295 6880 2304
rect 6828 2261 6837 2295
rect 6837 2261 6871 2295
rect 6871 2261 6880 2295
rect 6828 2252 6880 2261
rect 7380 2295 7432 2304
rect 7380 2261 7389 2295
rect 7389 2261 7423 2295
rect 7423 2261 7432 2295
rect 7380 2252 7432 2261
rect 7840 2320 7892 2372
rect 8208 2388 8260 2440
rect 8392 2320 8444 2372
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 9864 2456 9916 2508
rect 10416 2456 10468 2508
rect 8668 2320 8720 2372
rect 9588 2320 9640 2372
rect 10140 2320 10192 2372
rect 10968 2456 11020 2508
rect 11980 2567 12032 2576
rect 11980 2533 11989 2567
rect 11989 2533 12023 2567
rect 12023 2533 12032 2567
rect 11980 2524 12032 2533
rect 12256 2567 12308 2576
rect 12256 2533 12265 2567
rect 12265 2533 12299 2567
rect 12299 2533 12308 2567
rect 12256 2524 12308 2533
rect 12532 2567 12584 2576
rect 12532 2533 12541 2567
rect 12541 2533 12575 2567
rect 12575 2533 12584 2567
rect 12532 2524 12584 2533
rect 13820 2592 13872 2644
rect 13912 2635 13964 2644
rect 13912 2601 13921 2635
rect 13921 2601 13955 2635
rect 13955 2601 13964 2635
rect 13912 2592 13964 2601
rect 14188 2592 14240 2644
rect 18144 2592 18196 2644
rect 10692 2320 10744 2372
rect 11060 2388 11112 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 11428 2388 11480 2440
rect 12808 2456 12860 2508
rect 11244 2320 11296 2372
rect 11888 2320 11940 2372
rect 7932 2295 7984 2304
rect 7932 2261 7941 2295
rect 7941 2261 7975 2295
rect 7975 2261 7984 2295
rect 7932 2252 7984 2261
rect 8116 2252 8168 2304
rect 10324 2252 10376 2304
rect 10508 2295 10560 2304
rect 10508 2261 10517 2295
rect 10517 2261 10551 2295
rect 10551 2261 10560 2295
rect 10508 2252 10560 2261
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 11336 2295 11388 2304
rect 11336 2261 11345 2295
rect 11345 2261 11379 2295
rect 11379 2261 11388 2295
rect 11336 2252 11388 2261
rect 12716 2388 12768 2440
rect 12440 2320 12492 2372
rect 13544 2388 13596 2440
rect 16948 2524 17000 2576
rect 17040 2524 17092 2576
rect 19616 2592 19668 2644
rect 13452 2320 13504 2372
rect 13820 2388 13872 2440
rect 14832 2388 14884 2440
rect 15016 2388 15068 2440
rect 15292 2388 15344 2440
rect 15568 2388 15620 2440
rect 15844 2388 15896 2440
rect 16120 2388 16172 2440
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 17316 2388 17368 2440
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 19156 2456 19208 2508
rect 19340 2524 19392 2576
rect 23664 2592 23716 2644
rect 24768 2592 24820 2644
rect 26240 2592 26292 2644
rect 26884 2592 26936 2644
rect 28172 2592 28224 2644
rect 29000 2592 29052 2644
rect 29644 2592 29696 2644
rect 31760 2635 31812 2644
rect 31760 2601 31769 2635
rect 31769 2601 31803 2635
rect 31803 2601 31812 2635
rect 31760 2592 31812 2601
rect 17960 2388 18012 2440
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 18328 2388 18380 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19708 2388 19760 2440
rect 19892 2388 19944 2440
rect 22284 2456 22336 2508
rect 20904 2388 20956 2440
rect 21180 2388 21232 2440
rect 21548 2388 21600 2440
rect 22376 2388 22428 2440
rect 23572 2524 23624 2576
rect 27436 2524 27488 2576
rect 28908 2524 28960 2576
rect 30932 2524 30984 2576
rect 33508 2592 33560 2644
rect 35348 2592 35400 2644
rect 33416 2524 33468 2576
rect 35808 2524 35860 2576
rect 36728 2635 36780 2644
rect 36728 2601 36737 2635
rect 36737 2601 36771 2635
rect 36771 2601 36780 2635
rect 36728 2592 36780 2601
rect 36912 2592 36964 2644
rect 37004 2592 37056 2644
rect 37648 2524 37700 2576
rect 40040 2592 40092 2644
rect 40132 2635 40184 2644
rect 40132 2601 40141 2635
rect 40141 2601 40175 2635
rect 40175 2601 40184 2635
rect 40132 2592 40184 2601
rect 40224 2592 40276 2644
rect 40500 2592 40552 2644
rect 41696 2592 41748 2644
rect 43168 2592 43220 2644
rect 23480 2388 23532 2440
rect 23940 2388 23992 2440
rect 24860 2388 24912 2440
rect 25688 2388 25740 2440
rect 26240 2388 26292 2440
rect 26792 2431 26844 2440
rect 26792 2397 26801 2431
rect 26801 2397 26835 2431
rect 26835 2397 26844 2431
rect 26792 2388 26844 2397
rect 27068 2431 27120 2440
rect 27068 2397 27077 2431
rect 27077 2397 27111 2431
rect 27111 2397 27120 2431
rect 27068 2388 27120 2397
rect 12348 2252 12400 2304
rect 12808 2295 12860 2304
rect 12808 2261 12817 2295
rect 12817 2261 12851 2295
rect 12851 2261 12860 2295
rect 12808 2252 12860 2261
rect 14464 2252 14516 2304
rect 14832 2252 14884 2304
rect 15016 2252 15068 2304
rect 15108 2295 15160 2304
rect 15108 2261 15117 2295
rect 15117 2261 15151 2295
rect 15151 2261 15160 2295
rect 15108 2252 15160 2261
rect 15200 2252 15252 2304
rect 15568 2252 15620 2304
rect 15844 2252 15896 2304
rect 16120 2252 16172 2304
rect 16580 2320 16632 2372
rect 16672 2252 16724 2304
rect 17316 2252 17368 2304
rect 19524 2320 19576 2372
rect 18144 2252 18196 2304
rect 20352 2320 20404 2372
rect 21456 2320 21508 2372
rect 21640 2363 21692 2372
rect 21640 2329 21649 2363
rect 21649 2329 21683 2363
rect 21683 2329 21692 2363
rect 21640 2320 21692 2329
rect 24400 2320 24452 2372
rect 20720 2252 20772 2304
rect 22284 2295 22336 2304
rect 22284 2261 22293 2295
rect 22293 2261 22327 2295
rect 22327 2261 22336 2295
rect 22284 2252 22336 2261
rect 22836 2295 22888 2304
rect 22836 2261 22845 2295
rect 22845 2261 22879 2295
rect 22879 2261 22888 2295
rect 22836 2252 22888 2261
rect 23572 2295 23624 2304
rect 23572 2261 23581 2295
rect 23581 2261 23615 2295
rect 23615 2261 23624 2295
rect 23572 2252 23624 2261
rect 23664 2252 23716 2304
rect 24032 2252 24084 2304
rect 24952 2320 25004 2372
rect 27896 2388 27948 2440
rect 28080 2388 28132 2440
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 29368 2431 29420 2440
rect 29368 2397 29377 2431
rect 29377 2397 29411 2431
rect 29411 2397 29420 2431
rect 29368 2388 29420 2397
rect 29552 2388 29604 2440
rect 29828 2388 29880 2440
rect 31116 2320 31168 2372
rect 34336 2456 34388 2508
rect 34152 2388 34204 2440
rect 35992 2388 36044 2440
rect 36084 2388 36136 2440
rect 36544 2431 36596 2440
rect 36544 2397 36553 2431
rect 36553 2397 36587 2431
rect 36587 2397 36596 2431
rect 36544 2388 36596 2397
rect 36820 2456 36872 2508
rect 36912 2388 36964 2440
rect 37004 2431 37056 2440
rect 37004 2397 37013 2431
rect 37013 2397 37047 2431
rect 37047 2397 37056 2431
rect 37004 2388 37056 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 32128 2320 32180 2372
rect 32220 2363 32272 2372
rect 32220 2329 32229 2363
rect 32229 2329 32263 2363
rect 32263 2329 32272 2363
rect 32220 2320 32272 2329
rect 32404 2320 32456 2372
rect 33324 2363 33376 2372
rect 33324 2329 33333 2363
rect 33333 2329 33367 2363
rect 33367 2329 33376 2363
rect 33324 2320 33376 2329
rect 33876 2363 33928 2372
rect 33876 2329 33885 2363
rect 33885 2329 33919 2363
rect 33919 2329 33928 2363
rect 33876 2320 33928 2329
rect 34796 2363 34848 2372
rect 34796 2329 34805 2363
rect 34805 2329 34839 2363
rect 34839 2329 34848 2363
rect 34796 2320 34848 2329
rect 35348 2363 35400 2372
rect 35348 2329 35357 2363
rect 35357 2329 35391 2363
rect 35391 2329 35400 2363
rect 35348 2320 35400 2329
rect 36452 2320 36504 2372
rect 38384 2431 38436 2440
rect 38384 2397 38393 2431
rect 38393 2397 38427 2431
rect 38427 2397 38436 2431
rect 38384 2388 38436 2397
rect 38660 2431 38712 2440
rect 38660 2397 38669 2431
rect 38669 2397 38703 2431
rect 38703 2397 38712 2431
rect 38660 2388 38712 2397
rect 39120 2388 39172 2440
rect 39672 2431 39724 2440
rect 39672 2397 39681 2431
rect 39681 2397 39715 2431
rect 39715 2397 39724 2431
rect 39672 2388 39724 2397
rect 39764 2388 39816 2440
rect 40316 2431 40368 2440
rect 40316 2397 40325 2431
rect 40325 2397 40359 2431
rect 40359 2397 40368 2431
rect 40316 2388 40368 2397
rect 40408 2388 40460 2440
rect 40868 2431 40920 2440
rect 40868 2397 40877 2431
rect 40877 2397 40911 2431
rect 40911 2397 40920 2431
rect 40868 2388 40920 2397
rect 25504 2252 25556 2304
rect 26332 2252 26384 2304
rect 28356 2252 28408 2304
rect 30196 2252 30248 2304
rect 31668 2252 31720 2304
rect 32864 2252 32916 2304
rect 34152 2252 34204 2304
rect 34980 2252 35032 2304
rect 37096 2252 37148 2304
rect 38476 2320 38528 2372
rect 37832 2252 37884 2304
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38568 2295 38620 2304
rect 38568 2261 38577 2295
rect 38577 2261 38611 2295
rect 38611 2261 38620 2295
rect 38568 2252 38620 2261
rect 38936 2252 38988 2304
rect 39948 2320 40000 2372
rect 11644 2150 11696 2202
rect 11708 2150 11760 2202
rect 11772 2150 11824 2202
rect 11836 2150 11888 2202
rect 11900 2150 11952 2202
rect 22338 2150 22390 2202
rect 22402 2150 22454 2202
rect 22466 2150 22518 2202
rect 22530 2150 22582 2202
rect 22594 2150 22646 2202
rect 33032 2150 33084 2202
rect 33096 2150 33148 2202
rect 33160 2150 33212 2202
rect 33224 2150 33276 2202
rect 33288 2150 33340 2202
rect 43726 2150 43778 2202
rect 43790 2150 43842 2202
rect 43854 2150 43906 2202
rect 43918 2150 43970 2202
rect 43982 2150 44034 2202
rect 4896 2048 4948 2100
rect 5540 2048 5592 2100
rect 5908 2048 5960 2100
rect 10876 2048 10928 2100
rect 11428 2048 11480 2100
rect 19432 2048 19484 2100
rect 20812 2048 20864 2100
rect 20996 2048 21048 2100
rect 32404 2048 32456 2100
rect 11060 1980 11112 2032
rect 7932 1912 7984 1964
rect 8300 1912 8352 1964
rect 15200 1980 15252 2032
rect 16948 1980 17000 2032
rect 11336 1912 11388 1964
rect 13820 1844 13872 1896
rect 17684 1844 17736 1896
rect 18052 1844 18104 1896
rect 26792 1980 26844 2032
rect 29368 1980 29420 2032
rect 30380 1980 30432 2032
rect 32220 1980 32272 2032
rect 38292 2048 38344 2100
rect 38476 2048 38528 2100
rect 38568 2048 38620 2100
rect 21548 1844 21600 1896
rect 12164 1708 12216 1760
rect 6552 1640 6604 1692
rect 7380 1640 7432 1692
rect 8208 1640 8260 1692
rect 21916 1776 21968 1828
rect 32128 1844 32180 1896
rect 23020 1776 23072 1828
rect 31392 1708 31444 1760
rect 34980 1708 35032 1760
rect 35072 1708 35124 1760
rect 37004 1708 37056 1760
rect 12808 1640 12860 1692
rect 26424 1640 26476 1692
rect 16672 1572 16724 1624
rect 19156 1572 19208 1624
rect 38292 1572 38344 1624
rect 39672 1572 39724 1624
rect 8576 1504 8628 1556
rect 9312 1504 9364 1556
rect 17132 1504 17184 1556
rect 23204 1504 23256 1556
rect 34428 1504 34480 1556
rect 36544 1504 36596 1556
rect 37464 1504 37516 1556
rect 38476 1504 38528 1556
rect 39764 1504 39816 1556
rect 23756 1436 23808 1488
rect 31852 1436 31904 1488
rect 32864 1436 32916 1488
rect 35624 1436 35676 1488
rect 38568 1436 38620 1488
rect 40316 1436 40368 1488
rect 5632 1368 5684 1420
rect 6276 1368 6328 1420
rect 6828 1368 6880 1420
rect 11152 1368 11204 1420
rect 11796 1368 11848 1420
rect 12716 1368 12768 1420
rect 13176 1368 13228 1420
rect 32404 1368 32456 1420
rect 34152 1368 34204 1420
rect 37096 1368 37148 1420
rect 38384 1368 38436 1420
rect 39672 1368 39724 1420
rect 40868 1368 40920 1420
rect 15108 1300 15160 1352
rect 35348 1300 35400 1352
rect 15568 1232 15620 1284
rect 33784 1232 33836 1284
rect 16120 1164 16172 1216
rect 33692 1164 33744 1216
rect 15844 1096 15896 1148
rect 32036 1096 32088 1148
rect 17500 1028 17552 1080
rect 33876 1028 33928 1080
rect 23848 960 23900 1012
rect 10876 892 10928 944
rect 20076 892 20128 944
<< metal2 >>
rect 1306 9840 1362 10000
rect 3422 9840 3478 10000
rect 3528 9846 3832 9874
rect 1320 7546 1348 9840
rect 3436 9738 3464 9840
rect 3528 9738 3556 9846
rect 3436 9710 3556 9738
rect 3804 7546 3832 9846
rect 5538 9840 5594 10000
rect 7654 9840 7710 10000
rect 9770 9840 9826 10000
rect 11886 9840 11942 10000
rect 11992 9846 12204 9874
rect 5552 7546 5580 9840
rect 7668 7546 7696 9840
rect 9784 7546 9812 9840
rect 11900 9738 11928 9840
rect 11992 9738 12020 9846
rect 11900 9710 12020 9738
rect 11644 7644 11952 7653
rect 11644 7642 11650 7644
rect 11706 7642 11730 7644
rect 11786 7642 11810 7644
rect 11866 7642 11890 7644
rect 11946 7642 11952 7644
rect 11706 7590 11708 7642
rect 11888 7590 11890 7642
rect 11644 7588 11650 7590
rect 11706 7588 11730 7590
rect 11786 7588 11810 7590
rect 11866 7588 11890 7590
rect 11946 7588 11952 7590
rect 11644 7579 11952 7588
rect 12176 7546 12204 9846
rect 14002 9840 14058 10000
rect 16118 9840 16174 10000
rect 16224 9846 16528 9874
rect 14016 7546 14044 9840
rect 16132 9738 16160 9840
rect 16224 9738 16252 9846
rect 16132 9710 16252 9738
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 14004 7540 14056 7546
rect 16500 7528 16528 9846
rect 18234 9840 18290 10000
rect 20350 9840 20406 10000
rect 20456 9846 20668 9874
rect 16580 7540 16632 7546
rect 16500 7500 16580 7528
rect 14004 7482 14056 7488
rect 16580 7482 16632 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 4080 6186 4108 7346
rect 5736 6254 5764 7346
rect 6297 7100 6605 7109
rect 6297 7098 6303 7100
rect 6359 7098 6383 7100
rect 6439 7098 6463 7100
rect 6519 7098 6543 7100
rect 6599 7098 6605 7100
rect 6359 7046 6361 7098
rect 6541 7046 6543 7098
rect 6297 7044 6303 7046
rect 6359 7044 6383 7046
rect 6439 7044 6463 7046
rect 6519 7044 6543 7046
rect 6599 7044 6605 7046
rect 6297 7035 6605 7044
rect 11644 6556 11952 6565
rect 11644 6554 11650 6556
rect 11706 6554 11730 6556
rect 11786 6554 11810 6556
rect 11866 6554 11890 6556
rect 11946 6554 11952 6556
rect 11706 6502 11708 6554
rect 11888 6502 11890 6554
rect 11644 6500 11650 6502
rect 11706 6500 11730 6502
rect 11786 6500 11810 6502
rect 11866 6500 11890 6502
rect 11946 6500 11952 6502
rect 11644 6491 11952 6500
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 6297 6012 6605 6021
rect 6297 6010 6303 6012
rect 6359 6010 6383 6012
rect 6439 6010 6463 6012
rect 6519 6010 6543 6012
rect 6599 6010 6605 6012
rect 6359 5958 6361 6010
rect 6541 5958 6543 6010
rect 6297 5956 6303 5958
rect 6359 5956 6383 5958
rect 6439 5956 6463 5958
rect 6519 5956 6543 5958
rect 6599 5956 6605 5958
rect 6297 5947 6605 5956
rect 11644 5468 11952 5477
rect 11644 5466 11650 5468
rect 11706 5466 11730 5468
rect 11786 5466 11810 5468
rect 11866 5466 11890 5468
rect 11946 5466 11952 5468
rect 11706 5414 11708 5466
rect 11888 5414 11890 5466
rect 11644 5412 11650 5414
rect 11706 5412 11730 5414
rect 11786 5412 11810 5414
rect 11866 5412 11890 5414
rect 11946 5412 11952 5414
rect 11644 5403 11952 5412
rect 6297 4924 6605 4933
rect 6297 4922 6303 4924
rect 6359 4922 6383 4924
rect 6439 4922 6463 4924
rect 6519 4922 6543 4924
rect 6599 4922 6605 4924
rect 6359 4870 6361 4922
rect 6541 4870 6543 4922
rect 6297 4868 6303 4870
rect 6359 4868 6383 4870
rect 6439 4868 6463 4870
rect 6519 4868 6543 4870
rect 6599 4868 6605 4870
rect 6297 4859 6605 4868
rect 9680 4752 9732 4758
rect 7930 4720 7986 4729
rect 7852 4678 7930 4706
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6196 2582 6224 4558
rect 6297 3836 6605 3845
rect 6297 3834 6303 3836
rect 6359 3834 6383 3836
rect 6439 3834 6463 3836
rect 6519 3834 6543 3836
rect 6599 3834 6605 3836
rect 6359 3782 6361 3834
rect 6541 3782 6543 3834
rect 6297 3780 6303 3782
rect 6359 3780 6383 3782
rect 6439 3780 6463 3782
rect 6519 3780 6543 3782
rect 6599 3780 6605 3782
rect 6297 3771 6605 3780
rect 6297 2748 6605 2757
rect 6297 2746 6303 2748
rect 6359 2746 6383 2748
rect 6439 2746 6463 2748
rect 6519 2746 6543 2748
rect 6599 2746 6605 2748
rect 6359 2694 6361 2746
rect 6541 2694 6543 2746
rect 6297 2692 6303 2694
rect 6359 2692 6383 2694
rect 6439 2692 6463 2694
rect 6519 2692 6543 2694
rect 6599 2692 6605 2694
rect 6297 2683 6605 2692
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5552 2394 5580 2450
rect 4988 2372 5040 2378
rect 5264 2372 5316 2378
rect 5040 2332 5212 2360
rect 4988 2314 5040 2320
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4908 2106 4936 2246
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 5184 160 5212 2332
rect 5552 2366 5764 2394
rect 5316 2332 5488 2360
rect 5264 2314 5316 2320
rect 5460 160 5488 2332
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5552 2106 5580 2246
rect 5540 2100 5592 2106
rect 5540 2042 5592 2048
rect 5644 1426 5672 2246
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 5736 160 5764 2366
rect 5828 1306 5856 2450
rect 5920 2106 5948 2518
rect 6288 2514 6408 2530
rect 6276 2508 6408 2514
rect 6328 2502 6408 2508
rect 6276 2450 6328 2456
rect 5908 2100 5960 2106
rect 5908 2042 5960 2048
rect 6276 1420 6328 1426
rect 6276 1362 6328 1368
rect 5828 1278 6040 1306
rect 6012 160 6040 1278
rect 6288 160 6316 1362
rect 5170 0 5226 160
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6380 82 6408 2502
rect 6564 2446 6592 2586
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6564 1698 6592 2246
rect 6552 1692 6604 1698
rect 6552 1634 6604 1640
rect 6748 1306 6776 2450
rect 7380 2440 7432 2446
rect 7656 2440 7708 2446
rect 7432 2400 7512 2428
rect 7380 2382 7432 2388
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6840 1426 6868 2246
rect 6828 1420 6880 1426
rect 6828 1362 6880 1368
rect 6748 1278 6868 1306
rect 6840 160 6868 1278
rect 6550 82 6606 160
rect 6380 54 6606 82
rect 6550 0 6606 54
rect 6826 0 6882 160
rect 7024 82 7052 2314
rect 7102 82 7158 160
rect 7024 54 7158 82
rect 7300 82 7328 2314
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7392 1698 7420 2246
rect 7380 1692 7432 1698
rect 7380 1634 7432 1640
rect 7378 82 7434 160
rect 7300 54 7434 82
rect 7484 82 7512 2400
rect 7708 2400 7788 2428
rect 7656 2382 7708 2388
rect 7654 82 7710 160
rect 7484 54 7710 82
rect 7760 82 7788 2400
rect 7852 2378 7880 4678
rect 9680 4694 9732 4700
rect 7930 4655 7986 4664
rect 8206 4584 8262 4593
rect 8128 4542 8206 4570
rect 7932 2440 7984 2446
rect 7984 2400 8064 2428
rect 7932 2382 7984 2388
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7944 1970 7972 2246
rect 7932 1964 7984 1970
rect 7932 1906 7984 1912
rect 7930 82 7986 160
rect 7760 54 7986 82
rect 8036 82 8064 2400
rect 8128 2310 8156 4542
rect 8206 4519 8262 4528
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8680 2650 8708 4422
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9324 3194 9352 3538
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 8758 3088 8814 3097
rect 8758 3023 8814 3032
rect 9128 3052 9180 3058
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8220 1698 8248 2382
rect 8312 1970 8340 2518
rect 8772 2514 8800 3023
rect 9128 2994 9180 3000
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8392 2372 8444 2378
rect 8444 2332 8524 2360
rect 8392 2314 8444 2320
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8208 1692 8260 1698
rect 8208 1634 8260 1640
rect 8496 160 8524 2332
rect 8588 1562 8616 2382
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8576 1556 8628 1562
rect 8576 1498 8628 1504
rect 8206 82 8262 160
rect 8036 54 8262 82
rect 7102 0 7158 54
rect 7378 0 7434 54
rect 7654 0 7710 54
rect 7930 0 7986 54
rect 8206 0 8262 54
rect 8482 0 8538 160
rect 8680 82 8708 2314
rect 8758 82 8814 160
rect 8680 54 8814 82
rect 8758 0 8814 54
rect 9034 82 9090 160
rect 9140 82 9168 2994
rect 9692 2802 9720 4694
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9232 2774 9720 2802
rect 9232 2650 9260 2774
rect 9968 2650 9996 3878
rect 10244 2650 10272 4626
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 11644 4380 11952 4389
rect 11644 4378 11650 4380
rect 11706 4378 11730 4380
rect 11786 4378 11810 4380
rect 11866 4378 11890 4380
rect 11946 4378 11952 4380
rect 11706 4326 11708 4378
rect 11888 4326 11890 4378
rect 11644 4324 11650 4326
rect 11706 4324 11730 4326
rect 11786 4324 11810 4326
rect 11866 4324 11890 4326
rect 11946 4324 11952 4326
rect 11644 4315 11952 4324
rect 13912 4208 13964 4214
rect 13832 4156 13912 4162
rect 13832 4150 13964 4156
rect 13832 4134 13952 4150
rect 11978 4040 12034 4049
rect 10324 4004 10376 4010
rect 11978 3975 12034 3984
rect 10324 3946 10376 3952
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9324 160 9352 1498
rect 9416 1465 9444 2586
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 9402 1456 9458 1465
rect 9402 1391 9458 1400
rect 9600 160 9628 2314
rect 9876 160 9904 2450
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 10152 160 10180 2314
rect 10336 2310 10364 3946
rect 11058 3632 11114 3641
rect 11058 3567 11114 3576
rect 11072 2650 11100 3567
rect 11644 3292 11952 3301
rect 11644 3290 11650 3292
rect 11706 3290 11730 3292
rect 11786 3290 11810 3292
rect 11866 3290 11890 3292
rect 11946 3290 11952 3292
rect 11706 3238 11708 3290
rect 11888 3238 11890 3290
rect 11644 3236 11650 3238
rect 11706 3236 11730 3238
rect 11786 3236 11810 3238
rect 11866 3236 11890 3238
rect 11946 3236 11952 3238
rect 11644 3227 11952 3236
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11992 2582 12020 3975
rect 12530 3496 12586 3505
rect 12530 3431 12586 3440
rect 12544 2582 12572 3431
rect 13832 3074 13860 4134
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 13924 3194 13952 4014
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13832 3046 13952 3074
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13832 2650 13860 2926
rect 13924 2650 13952 3046
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 11980 2576 12032 2582
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 11072 2502 11560 2530
rect 11980 2518 12032 2524
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10428 160 10456 2450
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10520 1601 10548 2246
rect 10506 1592 10562 1601
rect 10506 1527 10562 1536
rect 10704 160 10732 2314
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 1193 10824 2246
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10782 1184 10838 1193
rect 10782 1119 10838 1128
rect 10888 950 10916 2042
rect 10876 944 10928 950
rect 10876 886 10928 892
rect 10980 160 11008 2450
rect 11072 2446 11100 2502
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11058 2272 11114 2281
rect 11058 2207 11114 2216
rect 11072 2038 11100 2207
rect 11060 2032 11112 2038
rect 11060 1974 11112 1980
rect 11164 1426 11192 2382
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 11256 160 11284 2314
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11348 1970 11376 2246
rect 11440 2106 11468 2382
rect 11428 2100 11480 2106
rect 11428 2042 11480 2048
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11532 160 11560 2502
rect 11888 2372 11940 2378
rect 11940 2332 12112 2360
rect 11888 2314 11940 2320
rect 11644 2204 11952 2213
rect 11644 2202 11650 2204
rect 11706 2202 11730 2204
rect 11786 2202 11810 2204
rect 11866 2202 11890 2204
rect 11946 2202 11952 2204
rect 11706 2150 11708 2202
rect 11888 2150 11890 2202
rect 11644 2148 11650 2150
rect 11706 2148 11730 2150
rect 11786 2148 11810 2150
rect 11866 2148 11890 2150
rect 11946 2148 11952 2150
rect 11644 2139 11952 2148
rect 11796 1420 11848 1426
rect 11796 1362 11848 1368
rect 11808 160 11836 1362
rect 12084 160 12112 2332
rect 12268 2281 12296 2518
rect 12808 2508 12860 2514
rect 12860 2468 12940 2496
rect 12808 2450 12860 2456
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12440 2372 12492 2378
rect 12492 2332 12664 2360
rect 12440 2314 12492 2320
rect 12348 2304 12400 2310
rect 12254 2272 12310 2281
rect 12348 2246 12400 2252
rect 12254 2207 12310 2216
rect 12162 2136 12218 2145
rect 12162 2071 12218 2080
rect 12176 1766 12204 2071
rect 12164 1760 12216 1766
rect 12164 1702 12216 1708
rect 12360 160 12388 2246
rect 12636 160 12664 2332
rect 12728 1426 12756 2382
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12820 1698 12848 2246
rect 12808 1692 12860 1698
rect 12808 1634 12860 1640
rect 12716 1420 12768 1426
rect 12716 1362 12768 1368
rect 12912 160 12940 2468
rect 13280 1873 13308 2586
rect 13544 2440 13596 2446
rect 13820 2440 13872 2446
rect 13596 2400 13768 2428
rect 13544 2382 13596 2388
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 13266 1864 13322 1873
rect 13266 1799 13322 1808
rect 13176 1420 13228 1426
rect 13176 1362 13228 1368
rect 13188 160 13216 1362
rect 13464 160 13492 2314
rect 13740 160 13768 2400
rect 13820 2382 13872 2388
rect 13832 1902 13860 2382
rect 13820 1896 13872 1902
rect 13820 1838 13872 1844
rect 14016 160 14044 2994
rect 14108 2990 14136 4490
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14200 2650 14228 7346
rect 16776 5914 16804 7346
rect 18248 7206 18276 9840
rect 20364 9738 20392 9840
rect 20456 9738 20484 9846
rect 20364 9710 20484 9738
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19076 7410 19104 7686
rect 20640 7426 20668 9846
rect 22466 9840 22522 10000
rect 22572 9846 22876 9874
rect 22480 9738 22508 9840
rect 22572 9738 22600 9846
rect 22480 9710 22600 9738
rect 22192 7812 22244 7818
rect 22192 7754 22244 7760
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20720 7472 20772 7478
rect 20640 7420 20720 7426
rect 20640 7414 20772 7420
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 19064 7404 19116 7410
rect 20640 7398 20760 7414
rect 19064 7346 19116 7352
rect 18616 7206 18644 7346
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 16991 7100 17299 7109
rect 16991 7098 16997 7100
rect 17053 7098 17077 7100
rect 17133 7098 17157 7100
rect 17213 7098 17237 7100
rect 17293 7098 17299 7100
rect 17053 7046 17055 7098
rect 17235 7046 17237 7098
rect 16991 7044 16997 7046
rect 17053 7044 17077 7046
rect 17133 7044 17157 7046
rect 17213 7044 17237 7046
rect 17293 7044 17299 7046
rect 16991 7035 17299 7044
rect 17328 7002 17356 7142
rect 21100 7002 21128 7482
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 16991 6012 17299 6021
rect 16991 6010 16997 6012
rect 17053 6010 17077 6012
rect 17133 6010 17157 6012
rect 17213 6010 17237 6012
rect 17293 6010 17299 6012
rect 17053 5958 17055 6010
rect 17235 5958 17237 6010
rect 16991 5956 16997 5958
rect 17053 5956 17077 5958
rect 17133 5956 17157 5958
rect 17213 5956 17237 5958
rect 17293 5956 17299 5958
rect 16991 5947 17299 5956
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16488 5704 16540 5710
rect 16486 5672 16488 5681
rect 16540 5672 16542 5681
rect 16486 5607 16542 5616
rect 16991 4924 17299 4933
rect 16991 4922 16997 4924
rect 17053 4922 17077 4924
rect 17133 4922 17157 4924
rect 17213 4922 17237 4924
rect 17293 4922 17299 4924
rect 17053 4870 17055 4922
rect 17235 4870 17237 4922
rect 16991 4868 16997 4870
rect 17053 4868 17077 4870
rect 17133 4868 17157 4870
rect 17213 4868 17237 4870
rect 17293 4868 17299 4870
rect 16991 4859 17299 4868
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14384 2774 14412 2994
rect 14292 2746 14412 2774
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14292 160 14320 2746
rect 14476 2310 14504 4218
rect 16991 3836 17299 3845
rect 16991 3834 16997 3836
rect 17053 3834 17077 3836
rect 17133 3834 17157 3836
rect 17213 3834 17237 3836
rect 17293 3834 17299 3836
rect 17053 3782 17055 3834
rect 17235 3782 17237 3834
rect 16991 3780 16997 3782
rect 17053 3780 17077 3782
rect 17133 3780 17157 3782
rect 17213 3780 17237 3782
rect 17293 3780 17299 3782
rect 16991 3771 17299 3780
rect 19154 3768 19210 3777
rect 15108 3732 15160 3738
rect 19154 3703 19210 3712
rect 15108 3674 15160 3680
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 9034 54 9168 82
rect 9034 0 9090 54
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10138 0 10194 160
rect 10414 0 10470 160
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11242 0 11298 160
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 82 14610 160
rect 14660 82 14688 2994
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14844 2310 14872 2382
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 921 14872 2246
rect 14830 912 14886 921
rect 14830 847 14886 856
rect 14554 54 14688 82
rect 14830 82 14886 160
rect 14936 82 14964 2994
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 15028 2446 15056 2858
rect 15120 2854 15148 3674
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15304 2446 15332 2790
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 14830 54 14964 82
rect 15028 82 15056 2246
rect 15120 1358 15148 2246
rect 15212 2038 15240 2246
rect 15200 2032 15252 2038
rect 15200 1974 15252 1980
rect 15108 1352 15160 1358
rect 15108 1294 15160 1300
rect 15396 160 15424 2994
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15580 2446 15608 2790
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15580 1290 15608 2246
rect 15568 1284 15620 1290
rect 15568 1226 15620 1232
rect 15672 160 15700 2994
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15856 2446 15884 2790
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15856 1154 15884 2246
rect 15844 1148 15896 1154
rect 15844 1090 15896 1096
rect 15948 160 15976 2994
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16132 2446 16160 2790
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16132 1222 16160 2246
rect 16120 1216 16172 1222
rect 16120 1158 16172 1164
rect 16224 160 16252 2994
rect 16316 2446 16344 3334
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16500 160 16528 2994
rect 16684 2446 16712 3606
rect 16764 3528 16816 3534
rect 17592 3528 17644 3534
rect 16764 3470 16816 3476
rect 17420 3488 17592 3516
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16592 1034 16620 2314
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16684 1630 16712 2246
rect 16672 1624 16724 1630
rect 16672 1566 16724 1572
rect 16670 1048 16726 1057
rect 16592 1006 16670 1034
rect 16670 983 16726 992
rect 16776 160 16804 3470
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16960 2938 16988 2994
rect 16868 2910 16988 2938
rect 16868 1578 16896 2910
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 16991 2748 17299 2757
rect 16991 2746 16997 2748
rect 17053 2746 17077 2748
rect 17133 2746 17157 2748
rect 17213 2746 17237 2748
rect 17293 2746 17299 2748
rect 17053 2694 17055 2746
rect 17235 2694 17237 2746
rect 16991 2692 16997 2694
rect 17053 2692 17077 2694
rect 17133 2692 17157 2694
rect 17213 2692 17237 2694
rect 17293 2692 17299 2694
rect 16991 2683 17299 2692
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 17040 2576 17092 2582
rect 17092 2524 17172 2530
rect 17040 2518 17172 2524
rect 16960 2038 16988 2518
rect 17052 2502 17172 2518
rect 16948 2032 17000 2038
rect 16948 1974 17000 1980
rect 16868 1550 17080 1578
rect 17144 1562 17172 2502
rect 17328 2446 17356 2790
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 1737 17356 2246
rect 17314 1728 17370 1737
rect 17314 1663 17370 1672
rect 17052 160 17080 1550
rect 17132 1556 17184 1562
rect 17132 1498 17184 1504
rect 15106 82 15162 160
rect 15028 54 15162 82
rect 14554 0 14610 54
rect 14830 0 14886 54
rect 15106 0 15162 54
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 0 16266 160
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 82 17370 160
rect 17420 82 17448 3488
rect 17592 3470 17644 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 17776 3392 17828 3398
rect 17696 3352 17776 3380
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17512 2938 17540 2994
rect 17512 2910 17632 2938
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17512 1086 17540 2790
rect 17500 1080 17552 1086
rect 17500 1022 17552 1028
rect 17604 160 17632 2910
rect 17696 2774 17724 3352
rect 17776 3334 17828 3340
rect 18234 3224 18290 3233
rect 18234 3159 18290 3168
rect 18052 3120 18104 3126
rect 18052 3062 18104 3068
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17788 2836 17816 2994
rect 17788 2808 17908 2836
rect 17696 2746 17816 2774
rect 17788 2446 17816 2746
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17696 1902 17724 2382
rect 17684 1896 17736 1902
rect 17684 1838 17736 1844
rect 17880 160 17908 2808
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 17972 1204 18000 2382
rect 18064 1902 18092 3062
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18156 2650 18184 2994
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18248 2530 18276 3159
rect 18326 2952 18382 2961
rect 18326 2887 18328 2896
rect 18380 2887 18382 2896
rect 18328 2858 18380 2864
rect 18156 2502 18276 2530
rect 18156 2310 18184 2502
rect 18236 2440 18288 2446
rect 18234 2408 18236 2417
rect 18328 2440 18380 2446
rect 18288 2408 18290 2417
rect 18328 2382 18380 2388
rect 18234 2343 18290 2352
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 18340 2145 18368 2382
rect 18326 2136 18382 2145
rect 18326 2071 18382 2080
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 17972 1176 18184 1204
rect 18156 160 18184 1176
rect 18432 160 18460 3470
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18616 3210 18644 3402
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18524 3182 18644 3210
rect 18524 1850 18552 3182
rect 18800 3058 18828 3334
rect 19168 3194 19196 3703
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18616 1986 18644 2994
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18892 2553 18920 2790
rect 18878 2544 18934 2553
rect 18878 2479 18934 2488
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19168 2009 19196 2450
rect 19154 2000 19210 2009
rect 18616 1958 19012 1986
rect 18524 1822 18736 1850
rect 18708 160 18736 1822
rect 18984 160 19012 1958
rect 19154 1935 19210 1944
rect 19156 1624 19208 1630
rect 19156 1566 19208 1572
rect 19168 1329 19196 1566
rect 19154 1320 19210 1329
rect 19154 1255 19210 1264
rect 19260 160 19288 3470
rect 19444 3466 19472 4694
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 20180 3534 20208 3878
rect 21744 3534 21772 3878
rect 19892 3528 19944 3534
rect 20168 3528 20220 3534
rect 19944 3488 20116 3516
rect 19892 3470 19944 3476
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19352 3194 19380 3334
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19616 3052 19668 3058
rect 19616 2994 19668 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19352 2582 19380 2926
rect 19628 2650 19656 2994
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 19720 2446 19748 3334
rect 19996 3194 20024 3334
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 19800 2916 19852 2922
rect 19800 2858 19852 2864
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 19444 2106 19472 2382
rect 19524 2372 19576 2378
rect 19524 2314 19576 2320
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19536 160 19564 2314
rect 19812 160 19840 2858
rect 19904 2446 19932 2994
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 20088 950 20116 3488
rect 20168 3470 20220 3476
rect 20812 3528 20864 3534
rect 21364 3528 21416 3534
rect 20864 3488 21128 3516
rect 20812 3470 20864 3476
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20824 3194 20852 3334
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20076 944 20128 950
rect 20076 886 20128 892
rect 17314 54 17448 82
rect 17314 0 17370 54
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 0 19026 160
rect 19246 0 19302 160
rect 19522 0 19578 160
rect 19798 0 19854 160
rect 20074 82 20130 160
rect 20272 82 20300 2790
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 20364 160 20392 2314
rect 20640 160 20668 2790
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 20074 54 20300 82
rect 20074 0 20130 54
rect 20350 0 20406 160
rect 20626 0 20682 160
rect 20732 82 20760 2246
rect 20824 2106 20852 2994
rect 20916 2446 20944 3334
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 21008 2106 21036 2858
rect 20812 2100 20864 2106
rect 20812 2042 20864 2048
rect 20996 2100 21048 2106
rect 20996 2042 21048 2048
rect 21100 1465 21128 3488
rect 21364 3470 21416 3476
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21192 2446 21220 3334
rect 21376 3097 21404 3470
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21468 3194 21496 3334
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21362 3088 21418 3097
rect 21362 3023 21418 3032
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21086 1456 21142 1465
rect 21086 1391 21142 1400
rect 20902 82 20958 160
rect 20732 54 20958 82
rect 20902 0 20958 54
rect 21178 82 21234 160
rect 21376 82 21404 2790
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 21468 160 21496 2314
rect 21560 1902 21588 2382
rect 21640 2372 21692 2378
rect 21640 2314 21692 2320
rect 21548 1896 21600 1902
rect 21548 1838 21600 1844
rect 21178 54 21404 82
rect 21178 0 21234 54
rect 21454 0 21510 160
rect 21652 82 21680 2314
rect 21928 1834 21956 7346
rect 22204 7274 22232 7754
rect 22338 7644 22646 7653
rect 22338 7642 22344 7644
rect 22400 7642 22424 7644
rect 22480 7642 22504 7644
rect 22560 7642 22584 7644
rect 22640 7642 22646 7644
rect 22400 7590 22402 7642
rect 22582 7590 22584 7642
rect 22338 7588 22344 7590
rect 22400 7588 22424 7590
rect 22480 7588 22504 7590
rect 22560 7588 22584 7590
rect 22640 7588 22646 7590
rect 22338 7579 22646 7588
rect 22848 7546 22876 9846
rect 24582 9840 24638 10000
rect 26698 9840 26754 10000
rect 28814 9840 28870 10000
rect 30930 9840 30986 10000
rect 33046 9840 33102 10000
rect 35162 9840 35218 10000
rect 37278 9840 37334 10000
rect 39394 9840 39450 10000
rect 39500 9846 39712 9874
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 24596 7426 24624 9840
rect 26712 7546 26740 9840
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 24688 7426 24716 7482
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23480 7404 23532 7410
rect 24596 7398 24716 7426
rect 28828 7426 28856 9840
rect 30944 7546 30972 9840
rect 33060 8514 33088 9840
rect 32968 8486 33088 8514
rect 31392 7812 31444 7818
rect 31392 7754 31444 7760
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 28920 7426 28948 7482
rect 24860 7404 24912 7410
rect 23480 7346 23532 7352
rect 24860 7346 24912 7352
rect 26884 7404 26936 7410
rect 28828 7398 28948 7426
rect 29000 7404 29052 7410
rect 26884 7346 26936 7352
rect 29000 7346 29052 7352
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 23400 7002 23428 7346
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23492 6798 23520 7346
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 22338 6556 22646 6565
rect 22338 6554 22344 6556
rect 22400 6554 22424 6556
rect 22480 6554 22504 6556
rect 22560 6554 22584 6556
rect 22640 6554 22646 6556
rect 22400 6502 22402 6554
rect 22582 6502 22584 6554
rect 22338 6500 22344 6502
rect 22400 6500 22424 6502
rect 22480 6500 22504 6502
rect 22560 6500 22584 6502
rect 22640 6500 22646 6502
rect 22338 6491 22646 6500
rect 22338 5468 22646 5477
rect 22338 5466 22344 5468
rect 22400 5466 22424 5468
rect 22480 5466 22504 5468
rect 22560 5466 22584 5468
rect 22640 5466 22646 5468
rect 22400 5414 22402 5466
rect 22582 5414 22584 5466
rect 22338 5412 22344 5414
rect 22400 5412 22424 5414
rect 22480 5412 22504 5414
rect 22560 5412 22584 5414
rect 22640 5412 22646 5414
rect 22338 5403 22646 5412
rect 22098 4720 22154 4729
rect 22098 4655 22154 4664
rect 22006 4584 22062 4593
rect 22006 4519 22062 4528
rect 22020 3534 22048 4519
rect 22112 3602 22140 4655
rect 22338 4380 22646 4389
rect 22338 4378 22344 4380
rect 22400 4378 22424 4380
rect 22480 4378 22504 4380
rect 22560 4378 22584 4380
rect 22640 4378 22646 4380
rect 22400 4326 22402 4378
rect 22582 4326 22584 4378
rect 22338 4324 22344 4326
rect 22400 4324 22424 4326
rect 22480 4324 22504 4326
rect 22560 4324 22584 4326
rect 22640 4324 22646 4326
rect 22338 4315 22646 4324
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22928 3392 22980 3398
rect 22928 3334 22980 3340
rect 22020 3194 22048 3334
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 21916 1828 21968 1834
rect 21916 1770 21968 1776
rect 22020 160 22048 2858
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22112 2632 22140 2790
rect 22204 2774 22232 3334
rect 22338 3292 22646 3301
rect 22338 3290 22344 3292
rect 22400 3290 22424 3292
rect 22480 3290 22504 3292
rect 22560 3290 22584 3292
rect 22640 3290 22646 3292
rect 22400 3238 22402 3290
rect 22582 3238 22584 3290
rect 22338 3236 22344 3238
rect 22400 3236 22424 3238
rect 22480 3236 22504 3238
rect 22560 3236 22584 3238
rect 22640 3236 22646 3238
rect 22338 3227 22646 3236
rect 22940 3194 22968 3334
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 22836 2848 22888 2854
rect 22756 2796 22836 2802
rect 22756 2790 22888 2796
rect 22756 2774 22876 2790
rect 22204 2746 22416 2774
rect 22112 2604 22324 2632
rect 22296 2514 22324 2604
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22388 2446 22416 2746
rect 22376 2440 22428 2446
rect 22204 2366 22324 2394
rect 22376 2382 22428 2388
rect 21730 82 21786 160
rect 21652 54 21786 82
rect 21730 0 21786 54
rect 22006 0 22062 160
rect 22204 82 22232 2366
rect 22296 2310 22324 2366
rect 22284 2304 22336 2310
rect 22284 2246 22336 2252
rect 22338 2204 22646 2213
rect 22338 2202 22344 2204
rect 22400 2202 22424 2204
rect 22480 2202 22504 2204
rect 22560 2202 22584 2204
rect 22640 2202 22646 2204
rect 22400 2150 22402 2202
rect 22582 2150 22584 2202
rect 22338 2148 22344 2150
rect 22400 2148 22424 2150
rect 22480 2148 22504 2150
rect 22560 2148 22584 2150
rect 22640 2148 22646 2150
rect 22338 2139 22646 2148
rect 22282 82 22338 160
rect 22204 54 22338 82
rect 22282 0 22338 54
rect 22558 82 22614 160
rect 22756 82 22784 2774
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 22848 160 22876 2246
rect 23032 1834 23060 6734
rect 24872 5914 24900 7346
rect 26896 6934 26924 7346
rect 27685 7100 27993 7109
rect 27685 7098 27691 7100
rect 27747 7098 27771 7100
rect 27827 7098 27851 7100
rect 27907 7098 27931 7100
rect 27987 7098 27993 7100
rect 27747 7046 27749 7098
rect 27929 7046 27931 7098
rect 27685 7044 27691 7046
rect 27747 7044 27771 7046
rect 27827 7044 27851 7046
rect 27907 7044 27931 7046
rect 27987 7044 27993 7046
rect 27685 7035 27993 7044
rect 26884 6928 26936 6934
rect 26884 6870 26936 6876
rect 27685 6012 27993 6021
rect 27685 6010 27691 6012
rect 27747 6010 27771 6012
rect 27827 6010 27851 6012
rect 27907 6010 27931 6012
rect 27987 6010 27993 6012
rect 27747 5958 27749 6010
rect 27929 5958 27931 6010
rect 27685 5956 27691 5958
rect 27747 5956 27771 5958
rect 27827 5956 27851 5958
rect 27907 5956 27931 5958
rect 27987 5956 27993 5958
rect 27685 5947 27993 5956
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 27685 4924 27993 4933
rect 27685 4922 27691 4924
rect 27747 4922 27771 4924
rect 27827 4922 27851 4924
rect 27907 4922 27931 4924
rect 27987 4922 27993 4924
rect 27747 4870 27749 4922
rect 27929 4870 27931 4922
rect 27685 4868 27691 4870
rect 27747 4868 27771 4870
rect 27827 4868 27851 4870
rect 27907 4868 27931 4870
rect 27987 4868 27993 4870
rect 27685 4859 27993 4868
rect 28816 4684 28868 4690
rect 28816 4626 28868 4632
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 23480 3664 23532 3670
rect 23480 3606 23532 3612
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23020 1828 23072 1834
rect 23020 1770 23072 1776
rect 23124 160 23152 2790
rect 23216 1562 23244 3470
rect 23492 2446 23520 3606
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23664 3460 23716 3466
rect 23664 3402 23716 3408
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23584 2582 23612 2926
rect 23676 2650 23704 3402
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23572 2576 23624 2582
rect 23572 2518 23624 2524
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23572 2304 23624 2310
rect 23572 2246 23624 2252
rect 23664 2304 23716 2310
rect 23664 2246 23716 2252
rect 23204 1556 23256 1562
rect 23204 1498 23256 1504
rect 23584 1442 23612 2246
rect 23400 1414 23612 1442
rect 23400 160 23428 1414
rect 23676 160 23704 2246
rect 23768 1494 23796 2994
rect 23756 1488 23808 1494
rect 23756 1430 23808 1436
rect 23860 1018 23888 3470
rect 23940 3392 23992 3398
rect 23992 3352 24072 3380
rect 23940 3334 23992 3340
rect 24044 2774 24072 3352
rect 24228 3058 24256 4558
rect 25964 4548 26016 4554
rect 25964 4490 26016 4496
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24412 3126 24440 3334
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 24504 3058 24532 4422
rect 25504 4276 25556 4282
rect 25504 4218 25556 4224
rect 24950 4040 25006 4049
rect 24950 3975 25006 3984
rect 24964 3602 24992 3975
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 25424 3534 25452 3878
rect 25516 3534 25544 4218
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25412 3528 25464 3534
rect 25412 3470 25464 3476
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 25240 3194 25268 3334
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24492 2848 24544 2854
rect 24492 2790 24544 2796
rect 23952 2746 24072 2774
rect 23952 2446 23980 2746
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 24400 2372 24452 2378
rect 24400 2314 24452 2320
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 24044 1170 24072 2246
rect 23952 1142 24072 1170
rect 23848 1012 23900 1018
rect 23848 954 23900 960
rect 23952 160 23980 1142
rect 22558 54 22784 82
rect 22558 0 22614 54
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 82 24270 160
rect 24412 82 24440 2314
rect 24504 160 24532 2790
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24780 160 24808 2586
rect 24872 2446 24900 2926
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24964 2378 24992 2858
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 25596 2848 25648 2854
rect 25596 2790 25648 2796
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 25056 160 25084 2790
rect 25504 2304 25556 2310
rect 25504 2246 25556 2252
rect 24214 54 24440 82
rect 24214 0 24270 54
rect 24490 0 24546 160
rect 24766 0 24822 160
rect 25042 0 25098 160
rect 25318 82 25374 160
rect 25516 82 25544 2246
rect 25608 160 25636 2790
rect 25700 2446 25728 3606
rect 25976 3534 26004 4490
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 26252 3777 26280 3878
rect 27685 3836 27993 3845
rect 27685 3834 27691 3836
rect 27747 3834 27771 3836
rect 27827 3834 27851 3836
rect 27907 3834 27931 3836
rect 27987 3834 27993 3836
rect 27747 3782 27749 3834
rect 27929 3782 27931 3834
rect 27685 3780 27691 3782
rect 27747 3780 27771 3782
rect 27827 3780 27851 3782
rect 27907 3780 27931 3782
rect 27987 3780 27993 3782
rect 26238 3768 26294 3777
rect 27685 3771 27993 3780
rect 26238 3703 26294 3712
rect 27068 3732 27120 3738
rect 27068 3674 27120 3680
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 26240 3528 26292 3534
rect 26516 3528 26568 3534
rect 26292 3488 26464 3516
rect 26240 3470 26292 3476
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 25318 54 25544 82
rect 25318 0 25374 54
rect 25594 0 25650 160
rect 25870 82 25926 160
rect 26068 82 26096 2790
rect 26160 2428 26188 3334
rect 26344 3194 26372 3334
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 26252 2650 26280 2994
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 26240 2440 26292 2446
rect 26160 2400 26240 2428
rect 26240 2382 26292 2388
rect 26332 2304 26384 2310
rect 26332 2246 26384 2252
rect 26344 1442 26372 2246
rect 26436 1698 26464 3488
rect 26514 3496 26516 3505
rect 26792 3528 26844 3534
rect 26568 3496 26570 3505
rect 26792 3470 26844 3476
rect 26514 3431 26570 3440
rect 26700 3460 26752 3466
rect 26700 3402 26752 3408
rect 26712 3126 26740 3402
rect 26700 3120 26752 3126
rect 26700 3062 26752 3068
rect 26608 2848 26660 2854
rect 26804 2825 26832 3470
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 26896 3126 26924 3334
rect 26884 3120 26936 3126
rect 26884 3062 26936 3068
rect 26976 2916 27028 2922
rect 26976 2858 27028 2864
rect 26608 2790 26660 2796
rect 26790 2816 26846 2825
rect 26424 1692 26476 1698
rect 26424 1634 26476 1640
rect 26160 1414 26372 1442
rect 26160 160 26188 1414
rect 25870 54 26096 82
rect 25870 0 25926 54
rect 26146 0 26202 160
rect 26422 82 26478 160
rect 26620 82 26648 2790
rect 26790 2751 26846 2760
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 26792 2440 26844 2446
rect 26792 2382 26844 2388
rect 26804 2038 26832 2382
rect 26792 2032 26844 2038
rect 26792 1974 26844 1980
rect 26422 54 26648 82
rect 26698 82 26754 160
rect 26896 82 26924 2586
rect 26988 160 27016 2858
rect 27080 2446 27108 3674
rect 27988 3664 28040 3670
rect 27618 3632 27674 3641
rect 27988 3606 28040 3612
rect 27618 3567 27674 3576
rect 27632 3534 27660 3567
rect 27160 3528 27212 3534
rect 27160 3470 27212 3476
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27172 2009 27200 3470
rect 28000 3074 28028 3606
rect 28828 3534 28856 4626
rect 29012 3738 29040 7346
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 29000 3732 29052 3738
rect 29000 3674 29052 3680
rect 29828 3664 29880 3670
rect 29828 3606 29880 3612
rect 29552 3596 29604 3602
rect 29552 3538 29604 3544
rect 28264 3528 28316 3534
rect 28540 3528 28592 3534
rect 28316 3488 28488 3516
rect 28264 3470 28316 3476
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 28092 3194 28120 3334
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 28000 3046 28120 3074
rect 27528 2916 27580 2922
rect 27528 2858 27580 2864
rect 27436 2576 27488 2582
rect 27436 2518 27488 2524
rect 27158 2000 27214 2009
rect 27158 1935 27214 1944
rect 26698 54 26924 82
rect 26422 0 26478 54
rect 26698 0 26754 54
rect 26974 0 27030 160
rect 27250 82 27306 160
rect 27448 82 27476 2518
rect 27540 160 27568 2858
rect 27685 2748 27993 2757
rect 27685 2746 27691 2748
rect 27747 2746 27771 2748
rect 27827 2746 27851 2748
rect 27907 2746 27931 2748
rect 27987 2746 27993 2748
rect 27747 2694 27749 2746
rect 27929 2694 27931 2746
rect 27685 2692 27691 2694
rect 27747 2692 27771 2694
rect 27827 2692 27851 2694
rect 27907 2692 27931 2694
rect 27987 2692 27993 2694
rect 27685 2683 27993 2692
rect 27894 2544 27950 2553
rect 27894 2479 27950 2488
rect 27908 2446 27936 2479
rect 28092 2446 28120 3046
rect 28356 2848 28408 2854
rect 28276 2796 28356 2802
rect 28276 2790 28408 2796
rect 28276 2774 28396 2790
rect 28172 2644 28224 2650
rect 28172 2586 28224 2592
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28184 218 28212 2586
rect 28000 190 28212 218
rect 27250 54 27476 82
rect 27250 0 27306 54
rect 27526 0 27582 160
rect 27802 82 27858 160
rect 28000 82 28028 190
rect 27802 54 28028 82
rect 28078 82 28134 160
rect 28276 82 28304 2774
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 28368 160 28396 2246
rect 28460 1193 28488 3488
rect 28540 3470 28592 3476
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28552 1601 28580 3470
rect 28724 3460 28776 3466
rect 28724 3402 28776 3408
rect 28632 3392 28684 3398
rect 28632 3334 28684 3340
rect 28644 3194 28672 3334
rect 28632 3188 28684 3194
rect 28632 3130 28684 3136
rect 28736 2446 28764 3402
rect 28998 3088 29054 3097
rect 28908 3052 28960 3058
rect 28998 3023 29000 3032
rect 28908 2994 28960 3000
rect 29052 3023 29054 3032
rect 29000 2994 29052 3000
rect 28920 2938 28948 2994
rect 29092 2984 29144 2990
rect 29090 2952 29092 2961
rect 29144 2952 29146 2961
rect 28920 2910 29040 2938
rect 28908 2848 28960 2854
rect 28828 2796 28908 2802
rect 28828 2790 28960 2796
rect 28828 2774 28948 2790
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 28538 1592 28594 1601
rect 28538 1527 28594 1536
rect 28446 1184 28502 1193
rect 28446 1119 28502 1128
rect 28078 54 28304 82
rect 27802 0 27858 54
rect 28078 0 28134 54
rect 28354 0 28410 160
rect 28630 82 28686 160
rect 28828 82 28856 2774
rect 29012 2650 29040 2910
rect 29090 2887 29146 2896
rect 29460 2848 29512 2854
rect 29196 2796 29460 2802
rect 29196 2790 29512 2796
rect 29196 2774 29500 2790
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 28920 160 28948 2518
rect 29196 160 29224 2774
rect 29564 2446 29592 3538
rect 29736 2916 29788 2922
rect 29736 2858 29788 2864
rect 29644 2644 29696 2650
rect 29644 2586 29696 2592
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29380 2038 29408 2382
rect 29368 2032 29420 2038
rect 29368 1974 29420 1980
rect 28630 54 28856 82
rect 28630 0 28686 54
rect 28906 0 28962 160
rect 29182 0 29238 160
rect 29458 82 29514 160
rect 29656 82 29684 2586
rect 29748 160 29776 2858
rect 29840 2446 29868 3606
rect 30024 3058 30052 3878
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 30288 2916 30340 2922
rect 30288 2858 30340 2864
rect 29828 2440 29880 2446
rect 29828 2382 29880 2388
rect 30196 2304 30248 2310
rect 30196 2246 30248 2252
rect 29458 54 29684 82
rect 29458 0 29514 54
rect 29734 0 29790 160
rect 30010 82 30066 160
rect 30208 82 30236 2246
rect 30300 160 30328 2858
rect 30380 2032 30432 2038
rect 30380 1974 30432 1980
rect 30392 1737 30420 1974
rect 30378 1728 30434 1737
rect 30378 1663 30434 1672
rect 30576 160 30604 3130
rect 30932 2576 30984 2582
rect 30932 2518 30984 2524
rect 30944 1306 30972 2518
rect 31116 2372 31168 2378
rect 31116 2314 31168 2320
rect 30852 1278 30972 1306
rect 30852 160 30880 1278
rect 31128 160 31156 2314
rect 31404 1766 31432 7754
rect 32968 7546 32996 8486
rect 33032 7644 33340 7653
rect 33032 7642 33038 7644
rect 33094 7642 33118 7644
rect 33174 7642 33198 7644
rect 33254 7642 33278 7644
rect 33334 7642 33340 7644
rect 33094 7590 33096 7642
rect 33276 7590 33278 7642
rect 33032 7588 33038 7590
rect 33094 7588 33118 7590
rect 33174 7588 33198 7590
rect 33254 7588 33278 7590
rect 33334 7588 33340 7590
rect 33032 7579 33340 7588
rect 35176 7546 35204 9840
rect 35900 7744 35952 7750
rect 35900 7686 35952 7692
rect 32956 7540 33008 7546
rect 32956 7482 33008 7488
rect 35164 7540 35216 7546
rect 35164 7482 35216 7488
rect 31760 7404 31812 7410
rect 31760 7346 31812 7352
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 31772 2650 31800 7346
rect 34336 7336 34388 7342
rect 34336 7278 34388 7284
rect 33032 6556 33340 6565
rect 33032 6554 33038 6556
rect 33094 6554 33118 6556
rect 33174 6554 33198 6556
rect 33254 6554 33278 6556
rect 33334 6554 33340 6556
rect 33094 6502 33096 6554
rect 33276 6502 33278 6554
rect 33032 6500 33038 6502
rect 33094 6500 33118 6502
rect 33174 6500 33198 6502
rect 33254 6500 33278 6502
rect 33334 6500 33340 6502
rect 33032 6491 33340 6500
rect 33600 6180 33652 6186
rect 33600 6122 33652 6128
rect 33032 5468 33340 5477
rect 33032 5466 33038 5468
rect 33094 5466 33118 5468
rect 33174 5466 33198 5468
rect 33254 5466 33278 5468
rect 33334 5466 33340 5468
rect 33094 5414 33096 5466
rect 33276 5414 33278 5466
rect 33032 5412 33038 5414
rect 33094 5412 33118 5414
rect 33174 5412 33198 5414
rect 33254 5412 33278 5414
rect 33334 5412 33340 5414
rect 33032 5403 33340 5412
rect 33032 4380 33340 4389
rect 33032 4378 33038 4380
rect 33094 4378 33118 4380
rect 33174 4378 33198 4380
rect 33254 4378 33278 4380
rect 33334 4378 33340 4380
rect 33094 4326 33096 4378
rect 33276 4326 33278 4378
rect 33032 4324 33038 4326
rect 33094 4324 33118 4326
rect 33174 4324 33198 4326
rect 33254 4324 33278 4326
rect 33334 4324 33340 4326
rect 33032 4315 33340 4324
rect 33416 4208 33468 4214
rect 33416 4150 33468 4156
rect 32036 3460 32088 3466
rect 32036 3402 32088 3408
rect 31944 2916 31996 2922
rect 31944 2858 31996 2864
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 31392 1760 31444 1766
rect 31392 1702 31444 1708
rect 31680 1578 31708 2246
rect 31588 1550 31708 1578
rect 30010 54 30236 82
rect 30010 0 30066 54
rect 30286 0 30342 160
rect 30562 0 30618 160
rect 30838 0 30894 160
rect 31114 0 31170 160
rect 31390 82 31446 160
rect 31588 82 31616 1550
rect 31852 1488 31904 1494
rect 31680 1436 31852 1442
rect 31680 1430 31904 1436
rect 31680 1414 31892 1430
rect 31680 160 31708 1414
rect 31956 160 31984 2858
rect 32048 1154 32076 3402
rect 32772 3392 32824 3398
rect 32772 3334 32824 3340
rect 32312 3052 32364 3058
rect 32312 2994 32364 3000
rect 32324 2854 32352 2994
rect 32496 2916 32548 2922
rect 32496 2858 32548 2864
rect 32312 2848 32364 2854
rect 32310 2816 32312 2825
rect 32364 2816 32366 2825
rect 32310 2751 32366 2760
rect 32128 2372 32180 2378
rect 32128 2314 32180 2320
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 32404 2372 32456 2378
rect 32404 2314 32456 2320
rect 32140 1902 32168 2314
rect 32232 2038 32260 2314
rect 32416 2106 32444 2314
rect 32404 2100 32456 2106
rect 32404 2042 32456 2048
rect 32220 2032 32272 2038
rect 32220 1974 32272 1980
rect 32128 1896 32180 1902
rect 32128 1838 32180 1844
rect 32404 1420 32456 1426
rect 32404 1362 32456 1368
rect 32036 1148 32088 1154
rect 32036 1090 32088 1096
rect 31390 54 31616 82
rect 31390 0 31446 54
rect 31666 0 31722 160
rect 31942 0 31998 160
rect 32218 82 32274 160
rect 32416 82 32444 1362
rect 32508 160 32536 2858
rect 32784 160 32812 3334
rect 33032 3292 33340 3301
rect 33032 3290 33038 3292
rect 33094 3290 33118 3292
rect 33174 3290 33198 3292
rect 33254 3290 33278 3292
rect 33334 3290 33340 3292
rect 33094 3238 33096 3290
rect 33276 3238 33278 3290
rect 33032 3236 33038 3238
rect 33094 3236 33118 3238
rect 33174 3236 33198 3238
rect 33254 3236 33278 3238
rect 33334 3236 33340 3238
rect 33032 3227 33340 3236
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 33060 2360 33088 3130
rect 33428 3126 33456 4150
rect 33612 3738 33640 6122
rect 33600 3732 33652 3738
rect 33600 3674 33652 3680
rect 33508 3460 33560 3466
rect 33508 3402 33560 3408
rect 33416 3120 33468 3126
rect 33416 3062 33468 3068
rect 33520 2650 33548 3402
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 33784 3052 33836 3058
rect 33784 2994 33836 3000
rect 33600 2916 33652 2922
rect 33600 2858 33652 2864
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 33416 2576 33468 2582
rect 33416 2518 33468 2524
rect 32968 2332 33088 2360
rect 33322 2408 33378 2417
rect 33322 2343 33324 2352
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 32876 1494 32904 2246
rect 32864 1488 32916 1494
rect 32864 1430 32916 1436
rect 32218 54 32444 82
rect 32218 0 32274 54
rect 32494 0 32550 160
rect 32770 0 32826 160
rect 32968 82 32996 2332
rect 33376 2343 33378 2352
rect 33324 2314 33376 2320
rect 33032 2204 33340 2213
rect 33032 2202 33038 2204
rect 33094 2202 33118 2204
rect 33174 2202 33198 2204
rect 33254 2202 33278 2204
rect 33334 2202 33340 2204
rect 33094 2150 33096 2202
rect 33276 2150 33278 2202
rect 33032 2148 33038 2150
rect 33094 2148 33118 2150
rect 33174 2148 33198 2150
rect 33254 2148 33278 2150
rect 33334 2148 33340 2150
rect 33032 2139 33340 2148
rect 33046 82 33102 160
rect 32968 54 33102 82
rect 33046 0 33102 54
rect 33322 82 33378 160
rect 33428 82 33456 2518
rect 33612 160 33640 2858
rect 33704 1222 33732 2994
rect 33796 1290 33824 2994
rect 34348 2514 34376 7278
rect 34428 6928 34480 6934
rect 35360 6914 35388 7346
rect 35532 7336 35584 7342
rect 35532 7278 35584 7284
rect 34480 6886 34560 6914
rect 35360 6886 35480 6914
rect 34428 6870 34480 6876
rect 34532 3194 34560 6886
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 34520 3188 34572 3194
rect 34520 3130 34572 3136
rect 34992 3126 35020 3334
rect 34980 3120 35032 3126
rect 34980 3062 35032 3068
rect 35256 3120 35308 3126
rect 35256 3062 35308 3068
rect 35452 3074 35480 6886
rect 35544 3194 35572 7278
rect 35808 6248 35860 6254
rect 35808 6190 35860 6196
rect 35532 3188 35584 3194
rect 35532 3130 35584 3136
rect 35624 3188 35676 3194
rect 35624 3130 35676 3136
rect 35636 3074 35664 3130
rect 34704 2984 34756 2990
rect 34704 2926 34756 2932
rect 34336 2508 34388 2514
rect 34336 2450 34388 2456
rect 34152 2440 34204 2446
rect 34072 2400 34152 2428
rect 33876 2372 33928 2378
rect 33876 2314 33928 2320
rect 33784 1284 33836 1290
rect 33784 1226 33836 1232
rect 33692 1216 33744 1222
rect 33692 1158 33744 1164
rect 33888 1086 33916 2314
rect 33876 1080 33928 1086
rect 33876 1022 33928 1028
rect 33322 54 33456 82
rect 33322 0 33378 54
rect 33598 0 33654 160
rect 33874 82 33930 160
rect 34072 82 34100 2400
rect 34152 2382 34204 2388
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 34164 1426 34192 2246
rect 34428 1556 34480 1562
rect 34428 1498 34480 1504
rect 34152 1420 34204 1426
rect 34152 1362 34204 1368
rect 34440 160 34468 1498
rect 34716 160 34744 2926
rect 34796 2372 34848 2378
rect 34796 2314 34848 2320
rect 34808 1057 34836 2314
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 34992 1766 35020 2246
rect 34980 1760 35032 1766
rect 34980 1702 35032 1708
rect 35072 1760 35124 1766
rect 35072 1702 35124 1708
rect 34794 1048 34850 1057
rect 34794 983 34850 992
rect 35084 898 35112 1702
rect 34992 870 35112 898
rect 34992 160 35020 870
rect 35268 160 35296 3062
rect 35348 3052 35400 3058
rect 35452 3046 35664 3074
rect 35348 2994 35400 3000
rect 35360 2650 35388 2994
rect 35716 2984 35768 2990
rect 35716 2926 35768 2932
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 35348 2372 35400 2378
rect 35348 2314 35400 2320
rect 35360 1358 35388 2314
rect 35624 1488 35676 1494
rect 35624 1430 35676 1436
rect 35348 1352 35400 1358
rect 35348 1294 35400 1300
rect 33874 54 34100 82
rect 33874 0 33930 54
rect 34150 0 34206 160
rect 34426 0 34482 160
rect 34702 0 34758 160
rect 34978 0 35034 160
rect 35254 0 35310 160
rect 35530 82 35586 160
rect 35636 82 35664 1430
rect 35728 218 35756 2926
rect 35820 2582 35848 6190
rect 35912 5574 35940 7686
rect 37292 7546 37320 9840
rect 39408 9738 39436 9840
rect 39500 9738 39528 9846
rect 39408 9710 39528 9738
rect 39684 7546 39712 9846
rect 41510 9840 41566 10000
rect 43626 9840 43682 10000
rect 41524 7546 41552 9840
rect 43640 7546 43668 9840
rect 43726 7644 44034 7653
rect 43726 7642 43732 7644
rect 43788 7642 43812 7644
rect 43868 7642 43892 7644
rect 43948 7642 43972 7644
rect 44028 7642 44034 7644
rect 43788 7590 43790 7642
rect 43970 7590 43972 7642
rect 43726 7588 43732 7590
rect 43788 7588 43812 7590
rect 43868 7588 43892 7590
rect 43948 7588 43972 7590
rect 44028 7588 44034 7590
rect 43726 7579 44034 7588
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 39672 7540 39724 7546
rect 39672 7482 39724 7488
rect 41512 7540 41564 7546
rect 41512 7482 41564 7488
rect 43628 7540 43680 7546
rect 43628 7482 43680 7488
rect 40224 7404 40276 7410
rect 40224 7346 40276 7352
rect 41696 7404 41748 7410
rect 41696 7346 41748 7352
rect 43168 7404 43220 7410
rect 43168 7346 43220 7352
rect 40040 7268 40092 7274
rect 40040 7210 40092 7216
rect 38379 7100 38687 7109
rect 38379 7098 38385 7100
rect 38441 7098 38465 7100
rect 38521 7098 38545 7100
rect 38601 7098 38625 7100
rect 38681 7098 38687 7100
rect 38441 7046 38443 7098
rect 38623 7046 38625 7098
rect 38379 7044 38385 7046
rect 38441 7044 38465 7046
rect 38521 7044 38545 7046
rect 38601 7044 38625 7046
rect 38681 7044 38687 7046
rect 38379 7035 38687 7044
rect 36728 6996 36780 7002
rect 36728 6938 36780 6944
rect 35900 5568 35952 5574
rect 35900 5510 35952 5516
rect 35992 2916 36044 2922
rect 35992 2858 36044 2864
rect 35808 2576 35860 2582
rect 35808 2518 35860 2524
rect 36004 2446 36032 2858
rect 36084 2848 36136 2854
rect 36360 2848 36412 2854
rect 36084 2790 36136 2796
rect 36358 2816 36360 2825
rect 36412 2816 36414 2825
rect 36096 2446 36124 2790
rect 36358 2751 36414 2760
rect 36740 2650 36768 6938
rect 38379 6012 38687 6021
rect 38379 6010 38385 6012
rect 38441 6010 38465 6012
rect 38521 6010 38545 6012
rect 38601 6010 38625 6012
rect 38681 6010 38687 6012
rect 38441 5958 38443 6010
rect 38623 5958 38625 6010
rect 38379 5956 38385 5958
rect 38441 5956 38465 5958
rect 38521 5956 38545 5958
rect 38601 5956 38625 5958
rect 38681 5956 38687 5958
rect 38379 5947 38687 5956
rect 38936 5704 38988 5710
rect 38936 5646 38988 5652
rect 38016 5568 38068 5574
rect 38016 5510 38068 5516
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 36832 3126 36860 3470
rect 36912 3392 36964 3398
rect 36912 3334 36964 3340
rect 36820 3120 36872 3126
rect 36820 3062 36872 3068
rect 36924 2650 36952 3334
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 37188 2848 37240 2854
rect 37188 2790 37240 2796
rect 36728 2644 36780 2650
rect 36728 2586 36780 2592
rect 36912 2644 36964 2650
rect 36912 2586 36964 2592
rect 37004 2644 37056 2650
rect 37004 2586 37056 2592
rect 37016 2530 37044 2586
rect 36820 2508 36872 2514
rect 36820 2450 36872 2456
rect 36924 2502 37044 2530
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36452 2372 36504 2378
rect 36188 2332 36452 2360
rect 36188 1306 36216 2332
rect 36452 2314 36504 2320
rect 36556 1562 36584 2382
rect 36544 1556 36596 1562
rect 36544 1498 36596 1504
rect 36096 1278 36216 1306
rect 35728 190 35848 218
rect 35820 160 35848 190
rect 36096 160 36124 1278
rect 36832 354 36860 2450
rect 36924 2446 36952 2502
rect 36912 2440 36964 2446
rect 36912 2382 36964 2388
rect 37004 2440 37056 2446
rect 37004 2382 37056 2388
rect 37016 1766 37044 2382
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 37004 1760 37056 1766
rect 37004 1702 37056 1708
rect 37108 1578 37136 2246
rect 36556 326 36860 354
rect 36924 1550 37136 1578
rect 35530 54 35664 82
rect 35530 0 35586 54
rect 35806 0 35862 160
rect 36082 0 36138 160
rect 36358 82 36414 160
rect 36556 82 36584 326
rect 36924 218 36952 1550
rect 37096 1420 37148 1426
rect 37096 1362 37148 1368
rect 36832 190 36952 218
rect 36358 54 36584 82
rect 36634 82 36690 160
rect 36832 82 36860 190
rect 36634 54 36860 82
rect 36910 82 36966 160
rect 37108 82 37136 1362
rect 37200 160 37228 2790
rect 37648 2576 37700 2582
rect 37568 2536 37648 2564
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 37476 1562 37504 2382
rect 37464 1556 37516 1562
rect 37464 1498 37516 1504
rect 37568 1306 37596 2536
rect 37648 2518 37700 2524
rect 37476 1278 37596 1306
rect 37476 160 37504 1278
rect 37752 160 37780 2994
rect 37830 2680 37886 2689
rect 37830 2615 37886 2624
rect 37844 2310 37872 2615
rect 38028 2310 38056 5510
rect 38379 4924 38687 4933
rect 38379 4922 38385 4924
rect 38441 4922 38465 4924
rect 38521 4922 38545 4924
rect 38601 4922 38625 4924
rect 38681 4922 38687 4924
rect 38441 4870 38443 4922
rect 38623 4870 38625 4922
rect 38379 4868 38385 4870
rect 38441 4868 38465 4870
rect 38521 4868 38545 4870
rect 38601 4868 38625 4870
rect 38681 4868 38687 4870
rect 38379 4859 38687 4868
rect 38379 3836 38687 3845
rect 38379 3834 38385 3836
rect 38441 3834 38465 3836
rect 38521 3834 38545 3836
rect 38601 3834 38625 3836
rect 38681 3834 38687 3836
rect 38441 3782 38443 3834
rect 38623 3782 38625 3834
rect 38379 3780 38385 3782
rect 38441 3780 38465 3782
rect 38521 3780 38545 3782
rect 38601 3780 38625 3782
rect 38681 3780 38687 3782
rect 38379 3771 38687 3780
rect 38844 3052 38896 3058
rect 38844 2994 38896 3000
rect 38752 2848 38804 2854
rect 38752 2790 38804 2796
rect 38379 2748 38687 2757
rect 38379 2746 38385 2748
rect 38441 2746 38465 2748
rect 38521 2746 38545 2748
rect 38601 2746 38625 2748
rect 38681 2746 38687 2748
rect 38441 2694 38443 2746
rect 38623 2694 38625 2746
rect 38379 2692 38385 2694
rect 38441 2692 38465 2694
rect 38521 2692 38545 2694
rect 38601 2692 38625 2694
rect 38681 2692 38687 2694
rect 38379 2683 38687 2692
rect 38764 2564 38792 2790
rect 38672 2536 38792 2564
rect 38672 2446 38700 2536
rect 38384 2440 38436 2446
rect 38384 2382 38436 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 37832 2304 37884 2310
rect 37832 2246 37884 2252
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 38304 2106 38332 2246
rect 38292 2100 38344 2106
rect 38292 2042 38344 2048
rect 38292 1624 38344 1630
rect 38292 1566 38344 1572
rect 38304 1408 38332 1566
rect 38396 1426 38424 2382
rect 38476 2372 38528 2378
rect 38476 2314 38528 2320
rect 38488 2106 38516 2314
rect 38568 2304 38620 2310
rect 38568 2246 38620 2252
rect 38580 2106 38608 2246
rect 38476 2100 38528 2106
rect 38476 2042 38528 2048
rect 38568 2100 38620 2106
rect 38568 2042 38620 2048
rect 38476 1556 38528 1562
rect 38476 1498 38528 1504
rect 38028 1380 38332 1408
rect 38384 1420 38436 1426
rect 38028 160 38056 1380
rect 38384 1362 38436 1368
rect 38488 1306 38516 1498
rect 38568 1488 38620 1494
rect 38568 1430 38620 1436
rect 38304 1278 38516 1306
rect 38304 160 38332 1278
rect 38580 160 38608 1430
rect 38856 160 38884 2994
rect 38948 2310 38976 5646
rect 39396 3052 39448 3058
rect 39396 2994 39448 3000
rect 39120 2848 39172 2854
rect 39120 2790 39172 2796
rect 39132 2446 39160 2790
rect 39120 2440 39172 2446
rect 39120 2382 39172 2388
rect 38936 2304 38988 2310
rect 38936 2246 38988 2252
rect 39408 1578 39436 2994
rect 40052 2650 40080 7210
rect 40132 2984 40184 2990
rect 40132 2926 40184 2932
rect 40144 2650 40172 2926
rect 40236 2650 40264 7346
rect 40500 7336 40552 7342
rect 40500 7278 40552 7284
rect 40408 2848 40460 2854
rect 40408 2790 40460 2796
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40132 2644 40184 2650
rect 40132 2586 40184 2592
rect 40224 2644 40276 2650
rect 40224 2586 40276 2592
rect 40420 2446 40448 2790
rect 40512 2650 40540 7278
rect 41708 2650 41736 7346
rect 43180 2650 43208 7346
rect 43726 6556 44034 6565
rect 43726 6554 43732 6556
rect 43788 6554 43812 6556
rect 43868 6554 43892 6556
rect 43948 6554 43972 6556
rect 44028 6554 44034 6556
rect 43788 6502 43790 6554
rect 43970 6502 43972 6554
rect 43726 6500 43732 6502
rect 43788 6500 43812 6502
rect 43868 6500 43892 6502
rect 43948 6500 43972 6502
rect 44028 6500 44034 6502
rect 43726 6491 44034 6500
rect 43726 5468 44034 5477
rect 43726 5466 43732 5468
rect 43788 5466 43812 5468
rect 43868 5466 43892 5468
rect 43948 5466 43972 5468
rect 44028 5466 44034 5468
rect 43788 5414 43790 5466
rect 43970 5414 43972 5466
rect 43726 5412 43732 5414
rect 43788 5412 43812 5414
rect 43868 5412 43892 5414
rect 43948 5412 43972 5414
rect 44028 5412 44034 5414
rect 43726 5403 44034 5412
rect 43726 4380 44034 4389
rect 43726 4378 43732 4380
rect 43788 4378 43812 4380
rect 43868 4378 43892 4380
rect 43948 4378 43972 4380
rect 44028 4378 44034 4380
rect 43788 4326 43790 4378
rect 43970 4326 43972 4378
rect 43726 4324 43732 4326
rect 43788 4324 43812 4326
rect 43868 4324 43892 4326
rect 43948 4324 43972 4326
rect 44028 4324 44034 4326
rect 43726 4315 44034 4324
rect 43726 3292 44034 3301
rect 43726 3290 43732 3292
rect 43788 3290 43812 3292
rect 43868 3290 43892 3292
rect 43948 3290 43972 3292
rect 44028 3290 44034 3292
rect 43788 3238 43790 3290
rect 43970 3238 43972 3290
rect 43726 3236 43732 3238
rect 43788 3236 43812 3238
rect 43868 3236 43892 3238
rect 43948 3236 43972 3238
rect 44028 3236 44034 3238
rect 43726 3227 44034 3236
rect 40500 2644 40552 2650
rect 40500 2586 40552 2592
rect 41696 2644 41748 2650
rect 41696 2586 41748 2592
rect 43168 2644 43220 2650
rect 43168 2586 43220 2592
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 39764 2440 39816 2446
rect 39764 2382 39816 2388
rect 40316 2440 40368 2446
rect 40316 2382 40368 2388
rect 40408 2440 40460 2446
rect 40408 2382 40460 2388
rect 40868 2440 40920 2446
rect 40868 2382 40920 2388
rect 39684 1630 39712 2382
rect 39132 1550 39436 1578
rect 39672 1624 39724 1630
rect 39672 1566 39724 1572
rect 39776 1562 39804 2382
rect 39948 2372 40000 2378
rect 39948 2314 40000 2320
rect 39764 1556 39816 1562
rect 39132 160 39160 1550
rect 39764 1498 39816 1504
rect 39672 1420 39724 1426
rect 39408 1380 39672 1408
rect 39408 160 39436 1380
rect 39672 1362 39724 1368
rect 39684 190 39804 218
rect 39684 160 39712 190
rect 36910 54 37136 82
rect 36358 0 36414 54
rect 36634 0 36690 54
rect 36910 0 36966 54
rect 37186 0 37242 160
rect 37462 0 37518 160
rect 37738 0 37794 160
rect 38014 0 38070 160
rect 38290 0 38346 160
rect 38566 0 38622 160
rect 38842 0 38898 160
rect 39118 0 39174 160
rect 39394 0 39450 160
rect 39670 0 39726 160
rect 39776 82 39804 190
rect 39960 82 39988 2314
rect 40328 1494 40356 2382
rect 40316 1488 40368 1494
rect 40316 1430 40368 1436
rect 40880 1426 40908 2382
rect 43726 2204 44034 2213
rect 43726 2202 43732 2204
rect 43788 2202 43812 2204
rect 43868 2202 43892 2204
rect 43948 2202 43972 2204
rect 44028 2202 44034 2204
rect 43788 2150 43790 2202
rect 43970 2150 43972 2202
rect 43726 2148 43732 2150
rect 43788 2148 43812 2150
rect 43868 2148 43892 2150
rect 43948 2148 43972 2150
rect 44028 2148 44034 2150
rect 43726 2139 44034 2148
rect 40868 1420 40920 1426
rect 40868 1362 40920 1368
rect 39776 54 39988 82
<< via2 >>
rect 11650 7642 11706 7644
rect 11730 7642 11786 7644
rect 11810 7642 11866 7644
rect 11890 7642 11946 7644
rect 11650 7590 11696 7642
rect 11696 7590 11706 7642
rect 11730 7590 11760 7642
rect 11760 7590 11772 7642
rect 11772 7590 11786 7642
rect 11810 7590 11824 7642
rect 11824 7590 11836 7642
rect 11836 7590 11866 7642
rect 11890 7590 11900 7642
rect 11900 7590 11946 7642
rect 11650 7588 11706 7590
rect 11730 7588 11786 7590
rect 11810 7588 11866 7590
rect 11890 7588 11946 7590
rect 6303 7098 6359 7100
rect 6383 7098 6439 7100
rect 6463 7098 6519 7100
rect 6543 7098 6599 7100
rect 6303 7046 6349 7098
rect 6349 7046 6359 7098
rect 6383 7046 6413 7098
rect 6413 7046 6425 7098
rect 6425 7046 6439 7098
rect 6463 7046 6477 7098
rect 6477 7046 6489 7098
rect 6489 7046 6519 7098
rect 6543 7046 6553 7098
rect 6553 7046 6599 7098
rect 6303 7044 6359 7046
rect 6383 7044 6439 7046
rect 6463 7044 6519 7046
rect 6543 7044 6599 7046
rect 11650 6554 11706 6556
rect 11730 6554 11786 6556
rect 11810 6554 11866 6556
rect 11890 6554 11946 6556
rect 11650 6502 11696 6554
rect 11696 6502 11706 6554
rect 11730 6502 11760 6554
rect 11760 6502 11772 6554
rect 11772 6502 11786 6554
rect 11810 6502 11824 6554
rect 11824 6502 11836 6554
rect 11836 6502 11866 6554
rect 11890 6502 11900 6554
rect 11900 6502 11946 6554
rect 11650 6500 11706 6502
rect 11730 6500 11786 6502
rect 11810 6500 11866 6502
rect 11890 6500 11946 6502
rect 6303 6010 6359 6012
rect 6383 6010 6439 6012
rect 6463 6010 6519 6012
rect 6543 6010 6599 6012
rect 6303 5958 6349 6010
rect 6349 5958 6359 6010
rect 6383 5958 6413 6010
rect 6413 5958 6425 6010
rect 6425 5958 6439 6010
rect 6463 5958 6477 6010
rect 6477 5958 6489 6010
rect 6489 5958 6519 6010
rect 6543 5958 6553 6010
rect 6553 5958 6599 6010
rect 6303 5956 6359 5958
rect 6383 5956 6439 5958
rect 6463 5956 6519 5958
rect 6543 5956 6599 5958
rect 11650 5466 11706 5468
rect 11730 5466 11786 5468
rect 11810 5466 11866 5468
rect 11890 5466 11946 5468
rect 11650 5414 11696 5466
rect 11696 5414 11706 5466
rect 11730 5414 11760 5466
rect 11760 5414 11772 5466
rect 11772 5414 11786 5466
rect 11810 5414 11824 5466
rect 11824 5414 11836 5466
rect 11836 5414 11866 5466
rect 11890 5414 11900 5466
rect 11900 5414 11946 5466
rect 11650 5412 11706 5414
rect 11730 5412 11786 5414
rect 11810 5412 11866 5414
rect 11890 5412 11946 5414
rect 6303 4922 6359 4924
rect 6383 4922 6439 4924
rect 6463 4922 6519 4924
rect 6543 4922 6599 4924
rect 6303 4870 6349 4922
rect 6349 4870 6359 4922
rect 6383 4870 6413 4922
rect 6413 4870 6425 4922
rect 6425 4870 6439 4922
rect 6463 4870 6477 4922
rect 6477 4870 6489 4922
rect 6489 4870 6519 4922
rect 6543 4870 6553 4922
rect 6553 4870 6599 4922
rect 6303 4868 6359 4870
rect 6383 4868 6439 4870
rect 6463 4868 6519 4870
rect 6543 4868 6599 4870
rect 6303 3834 6359 3836
rect 6383 3834 6439 3836
rect 6463 3834 6519 3836
rect 6543 3834 6599 3836
rect 6303 3782 6349 3834
rect 6349 3782 6359 3834
rect 6383 3782 6413 3834
rect 6413 3782 6425 3834
rect 6425 3782 6439 3834
rect 6463 3782 6477 3834
rect 6477 3782 6489 3834
rect 6489 3782 6519 3834
rect 6543 3782 6553 3834
rect 6553 3782 6599 3834
rect 6303 3780 6359 3782
rect 6383 3780 6439 3782
rect 6463 3780 6519 3782
rect 6543 3780 6599 3782
rect 6303 2746 6359 2748
rect 6383 2746 6439 2748
rect 6463 2746 6519 2748
rect 6543 2746 6599 2748
rect 6303 2694 6349 2746
rect 6349 2694 6359 2746
rect 6383 2694 6413 2746
rect 6413 2694 6425 2746
rect 6425 2694 6439 2746
rect 6463 2694 6477 2746
rect 6477 2694 6489 2746
rect 6489 2694 6519 2746
rect 6543 2694 6553 2746
rect 6553 2694 6599 2746
rect 6303 2692 6359 2694
rect 6383 2692 6439 2694
rect 6463 2692 6519 2694
rect 6543 2692 6599 2694
rect 7930 4664 7986 4720
rect 8206 4528 8262 4584
rect 8758 3032 8814 3088
rect 11650 4378 11706 4380
rect 11730 4378 11786 4380
rect 11810 4378 11866 4380
rect 11890 4378 11946 4380
rect 11650 4326 11696 4378
rect 11696 4326 11706 4378
rect 11730 4326 11760 4378
rect 11760 4326 11772 4378
rect 11772 4326 11786 4378
rect 11810 4326 11824 4378
rect 11824 4326 11836 4378
rect 11836 4326 11866 4378
rect 11890 4326 11900 4378
rect 11900 4326 11946 4378
rect 11650 4324 11706 4326
rect 11730 4324 11786 4326
rect 11810 4324 11866 4326
rect 11890 4324 11946 4326
rect 11978 3984 12034 4040
rect 9402 1400 9458 1456
rect 11058 3576 11114 3632
rect 11650 3290 11706 3292
rect 11730 3290 11786 3292
rect 11810 3290 11866 3292
rect 11890 3290 11946 3292
rect 11650 3238 11696 3290
rect 11696 3238 11706 3290
rect 11730 3238 11760 3290
rect 11760 3238 11772 3290
rect 11772 3238 11786 3290
rect 11810 3238 11824 3290
rect 11824 3238 11836 3290
rect 11836 3238 11866 3290
rect 11890 3238 11900 3290
rect 11900 3238 11946 3290
rect 11650 3236 11706 3238
rect 11730 3236 11786 3238
rect 11810 3236 11866 3238
rect 11890 3236 11946 3238
rect 12530 3440 12586 3496
rect 10506 1536 10562 1592
rect 10782 1128 10838 1184
rect 11058 2216 11114 2272
rect 11650 2202 11706 2204
rect 11730 2202 11786 2204
rect 11810 2202 11866 2204
rect 11890 2202 11946 2204
rect 11650 2150 11696 2202
rect 11696 2150 11706 2202
rect 11730 2150 11760 2202
rect 11760 2150 11772 2202
rect 11772 2150 11786 2202
rect 11810 2150 11824 2202
rect 11824 2150 11836 2202
rect 11836 2150 11866 2202
rect 11890 2150 11900 2202
rect 11900 2150 11946 2202
rect 11650 2148 11706 2150
rect 11730 2148 11786 2150
rect 11810 2148 11866 2150
rect 11890 2148 11946 2150
rect 12254 2216 12310 2272
rect 12162 2080 12218 2136
rect 13266 1808 13322 1864
rect 16997 7098 17053 7100
rect 17077 7098 17133 7100
rect 17157 7098 17213 7100
rect 17237 7098 17293 7100
rect 16997 7046 17043 7098
rect 17043 7046 17053 7098
rect 17077 7046 17107 7098
rect 17107 7046 17119 7098
rect 17119 7046 17133 7098
rect 17157 7046 17171 7098
rect 17171 7046 17183 7098
rect 17183 7046 17213 7098
rect 17237 7046 17247 7098
rect 17247 7046 17293 7098
rect 16997 7044 17053 7046
rect 17077 7044 17133 7046
rect 17157 7044 17213 7046
rect 17237 7044 17293 7046
rect 16997 6010 17053 6012
rect 17077 6010 17133 6012
rect 17157 6010 17213 6012
rect 17237 6010 17293 6012
rect 16997 5958 17043 6010
rect 17043 5958 17053 6010
rect 17077 5958 17107 6010
rect 17107 5958 17119 6010
rect 17119 5958 17133 6010
rect 17157 5958 17171 6010
rect 17171 5958 17183 6010
rect 17183 5958 17213 6010
rect 17237 5958 17247 6010
rect 17247 5958 17293 6010
rect 16997 5956 17053 5958
rect 17077 5956 17133 5958
rect 17157 5956 17213 5958
rect 17237 5956 17293 5958
rect 16486 5652 16488 5672
rect 16488 5652 16540 5672
rect 16540 5652 16542 5672
rect 16486 5616 16542 5652
rect 16997 4922 17053 4924
rect 17077 4922 17133 4924
rect 17157 4922 17213 4924
rect 17237 4922 17293 4924
rect 16997 4870 17043 4922
rect 17043 4870 17053 4922
rect 17077 4870 17107 4922
rect 17107 4870 17119 4922
rect 17119 4870 17133 4922
rect 17157 4870 17171 4922
rect 17171 4870 17183 4922
rect 17183 4870 17213 4922
rect 17237 4870 17247 4922
rect 17247 4870 17293 4922
rect 16997 4868 17053 4870
rect 17077 4868 17133 4870
rect 17157 4868 17213 4870
rect 17237 4868 17293 4870
rect 16997 3834 17053 3836
rect 17077 3834 17133 3836
rect 17157 3834 17213 3836
rect 17237 3834 17293 3836
rect 16997 3782 17043 3834
rect 17043 3782 17053 3834
rect 17077 3782 17107 3834
rect 17107 3782 17119 3834
rect 17119 3782 17133 3834
rect 17157 3782 17171 3834
rect 17171 3782 17183 3834
rect 17183 3782 17213 3834
rect 17237 3782 17247 3834
rect 17247 3782 17293 3834
rect 16997 3780 17053 3782
rect 17077 3780 17133 3782
rect 17157 3780 17213 3782
rect 17237 3780 17293 3782
rect 19154 3712 19210 3768
rect 14830 856 14886 912
rect 16670 992 16726 1048
rect 16997 2746 17053 2748
rect 17077 2746 17133 2748
rect 17157 2746 17213 2748
rect 17237 2746 17293 2748
rect 16997 2694 17043 2746
rect 17043 2694 17053 2746
rect 17077 2694 17107 2746
rect 17107 2694 17119 2746
rect 17119 2694 17133 2746
rect 17157 2694 17171 2746
rect 17171 2694 17183 2746
rect 17183 2694 17213 2746
rect 17237 2694 17247 2746
rect 17247 2694 17293 2746
rect 16997 2692 17053 2694
rect 17077 2692 17133 2694
rect 17157 2692 17213 2694
rect 17237 2692 17293 2694
rect 17314 1672 17370 1728
rect 18234 3168 18290 3224
rect 18326 2916 18382 2952
rect 18326 2896 18328 2916
rect 18328 2896 18380 2916
rect 18380 2896 18382 2916
rect 18234 2388 18236 2408
rect 18236 2388 18288 2408
rect 18288 2388 18290 2408
rect 18234 2352 18290 2388
rect 18326 2080 18382 2136
rect 18878 2488 18934 2544
rect 19154 1944 19210 2000
rect 19154 1264 19210 1320
rect 21362 3032 21418 3088
rect 21086 1400 21142 1456
rect 22344 7642 22400 7644
rect 22424 7642 22480 7644
rect 22504 7642 22560 7644
rect 22584 7642 22640 7644
rect 22344 7590 22390 7642
rect 22390 7590 22400 7642
rect 22424 7590 22454 7642
rect 22454 7590 22466 7642
rect 22466 7590 22480 7642
rect 22504 7590 22518 7642
rect 22518 7590 22530 7642
rect 22530 7590 22560 7642
rect 22584 7590 22594 7642
rect 22594 7590 22640 7642
rect 22344 7588 22400 7590
rect 22424 7588 22480 7590
rect 22504 7588 22560 7590
rect 22584 7588 22640 7590
rect 22344 6554 22400 6556
rect 22424 6554 22480 6556
rect 22504 6554 22560 6556
rect 22584 6554 22640 6556
rect 22344 6502 22390 6554
rect 22390 6502 22400 6554
rect 22424 6502 22454 6554
rect 22454 6502 22466 6554
rect 22466 6502 22480 6554
rect 22504 6502 22518 6554
rect 22518 6502 22530 6554
rect 22530 6502 22560 6554
rect 22584 6502 22594 6554
rect 22594 6502 22640 6554
rect 22344 6500 22400 6502
rect 22424 6500 22480 6502
rect 22504 6500 22560 6502
rect 22584 6500 22640 6502
rect 22344 5466 22400 5468
rect 22424 5466 22480 5468
rect 22504 5466 22560 5468
rect 22584 5466 22640 5468
rect 22344 5414 22390 5466
rect 22390 5414 22400 5466
rect 22424 5414 22454 5466
rect 22454 5414 22466 5466
rect 22466 5414 22480 5466
rect 22504 5414 22518 5466
rect 22518 5414 22530 5466
rect 22530 5414 22560 5466
rect 22584 5414 22594 5466
rect 22594 5414 22640 5466
rect 22344 5412 22400 5414
rect 22424 5412 22480 5414
rect 22504 5412 22560 5414
rect 22584 5412 22640 5414
rect 22098 4664 22154 4720
rect 22006 4528 22062 4584
rect 22344 4378 22400 4380
rect 22424 4378 22480 4380
rect 22504 4378 22560 4380
rect 22584 4378 22640 4380
rect 22344 4326 22390 4378
rect 22390 4326 22400 4378
rect 22424 4326 22454 4378
rect 22454 4326 22466 4378
rect 22466 4326 22480 4378
rect 22504 4326 22518 4378
rect 22518 4326 22530 4378
rect 22530 4326 22560 4378
rect 22584 4326 22594 4378
rect 22594 4326 22640 4378
rect 22344 4324 22400 4326
rect 22424 4324 22480 4326
rect 22504 4324 22560 4326
rect 22584 4324 22640 4326
rect 22344 3290 22400 3292
rect 22424 3290 22480 3292
rect 22504 3290 22560 3292
rect 22584 3290 22640 3292
rect 22344 3238 22390 3290
rect 22390 3238 22400 3290
rect 22424 3238 22454 3290
rect 22454 3238 22466 3290
rect 22466 3238 22480 3290
rect 22504 3238 22518 3290
rect 22518 3238 22530 3290
rect 22530 3238 22560 3290
rect 22584 3238 22594 3290
rect 22594 3238 22640 3290
rect 22344 3236 22400 3238
rect 22424 3236 22480 3238
rect 22504 3236 22560 3238
rect 22584 3236 22640 3238
rect 22344 2202 22400 2204
rect 22424 2202 22480 2204
rect 22504 2202 22560 2204
rect 22584 2202 22640 2204
rect 22344 2150 22390 2202
rect 22390 2150 22400 2202
rect 22424 2150 22454 2202
rect 22454 2150 22466 2202
rect 22466 2150 22480 2202
rect 22504 2150 22518 2202
rect 22518 2150 22530 2202
rect 22530 2150 22560 2202
rect 22584 2150 22594 2202
rect 22594 2150 22640 2202
rect 22344 2148 22400 2150
rect 22424 2148 22480 2150
rect 22504 2148 22560 2150
rect 22584 2148 22640 2150
rect 27691 7098 27747 7100
rect 27771 7098 27827 7100
rect 27851 7098 27907 7100
rect 27931 7098 27987 7100
rect 27691 7046 27737 7098
rect 27737 7046 27747 7098
rect 27771 7046 27801 7098
rect 27801 7046 27813 7098
rect 27813 7046 27827 7098
rect 27851 7046 27865 7098
rect 27865 7046 27877 7098
rect 27877 7046 27907 7098
rect 27931 7046 27941 7098
rect 27941 7046 27987 7098
rect 27691 7044 27747 7046
rect 27771 7044 27827 7046
rect 27851 7044 27907 7046
rect 27931 7044 27987 7046
rect 27691 6010 27747 6012
rect 27771 6010 27827 6012
rect 27851 6010 27907 6012
rect 27931 6010 27987 6012
rect 27691 5958 27737 6010
rect 27737 5958 27747 6010
rect 27771 5958 27801 6010
rect 27801 5958 27813 6010
rect 27813 5958 27827 6010
rect 27851 5958 27865 6010
rect 27865 5958 27877 6010
rect 27877 5958 27907 6010
rect 27931 5958 27941 6010
rect 27941 5958 27987 6010
rect 27691 5956 27747 5958
rect 27771 5956 27827 5958
rect 27851 5956 27907 5958
rect 27931 5956 27987 5958
rect 27691 4922 27747 4924
rect 27771 4922 27827 4924
rect 27851 4922 27907 4924
rect 27931 4922 27987 4924
rect 27691 4870 27737 4922
rect 27737 4870 27747 4922
rect 27771 4870 27801 4922
rect 27801 4870 27813 4922
rect 27813 4870 27827 4922
rect 27851 4870 27865 4922
rect 27865 4870 27877 4922
rect 27877 4870 27907 4922
rect 27931 4870 27941 4922
rect 27941 4870 27987 4922
rect 27691 4868 27747 4870
rect 27771 4868 27827 4870
rect 27851 4868 27907 4870
rect 27931 4868 27987 4870
rect 24950 3984 25006 4040
rect 27691 3834 27747 3836
rect 27771 3834 27827 3836
rect 27851 3834 27907 3836
rect 27931 3834 27987 3836
rect 27691 3782 27737 3834
rect 27737 3782 27747 3834
rect 27771 3782 27801 3834
rect 27801 3782 27813 3834
rect 27813 3782 27827 3834
rect 27851 3782 27865 3834
rect 27865 3782 27877 3834
rect 27877 3782 27907 3834
rect 27931 3782 27941 3834
rect 27941 3782 27987 3834
rect 27691 3780 27747 3782
rect 27771 3780 27827 3782
rect 27851 3780 27907 3782
rect 27931 3780 27987 3782
rect 26238 3712 26294 3768
rect 26514 3476 26516 3496
rect 26516 3476 26568 3496
rect 26568 3476 26570 3496
rect 26514 3440 26570 3476
rect 26790 2760 26846 2816
rect 27618 3576 27674 3632
rect 27158 1944 27214 2000
rect 27691 2746 27747 2748
rect 27771 2746 27827 2748
rect 27851 2746 27907 2748
rect 27931 2746 27987 2748
rect 27691 2694 27737 2746
rect 27737 2694 27747 2746
rect 27771 2694 27801 2746
rect 27801 2694 27813 2746
rect 27813 2694 27827 2746
rect 27851 2694 27865 2746
rect 27865 2694 27877 2746
rect 27877 2694 27907 2746
rect 27931 2694 27941 2746
rect 27941 2694 27987 2746
rect 27691 2692 27747 2694
rect 27771 2692 27827 2694
rect 27851 2692 27907 2694
rect 27931 2692 27987 2694
rect 27894 2488 27950 2544
rect 28998 3052 29054 3088
rect 28998 3032 29000 3052
rect 29000 3032 29052 3052
rect 29052 3032 29054 3052
rect 28538 1536 28594 1592
rect 28446 1128 28502 1184
rect 29090 2932 29092 2952
rect 29092 2932 29144 2952
rect 29144 2932 29146 2952
rect 29090 2896 29146 2932
rect 30378 1672 30434 1728
rect 33038 7642 33094 7644
rect 33118 7642 33174 7644
rect 33198 7642 33254 7644
rect 33278 7642 33334 7644
rect 33038 7590 33084 7642
rect 33084 7590 33094 7642
rect 33118 7590 33148 7642
rect 33148 7590 33160 7642
rect 33160 7590 33174 7642
rect 33198 7590 33212 7642
rect 33212 7590 33224 7642
rect 33224 7590 33254 7642
rect 33278 7590 33288 7642
rect 33288 7590 33334 7642
rect 33038 7588 33094 7590
rect 33118 7588 33174 7590
rect 33198 7588 33254 7590
rect 33278 7588 33334 7590
rect 33038 6554 33094 6556
rect 33118 6554 33174 6556
rect 33198 6554 33254 6556
rect 33278 6554 33334 6556
rect 33038 6502 33084 6554
rect 33084 6502 33094 6554
rect 33118 6502 33148 6554
rect 33148 6502 33160 6554
rect 33160 6502 33174 6554
rect 33198 6502 33212 6554
rect 33212 6502 33224 6554
rect 33224 6502 33254 6554
rect 33278 6502 33288 6554
rect 33288 6502 33334 6554
rect 33038 6500 33094 6502
rect 33118 6500 33174 6502
rect 33198 6500 33254 6502
rect 33278 6500 33334 6502
rect 33038 5466 33094 5468
rect 33118 5466 33174 5468
rect 33198 5466 33254 5468
rect 33278 5466 33334 5468
rect 33038 5414 33084 5466
rect 33084 5414 33094 5466
rect 33118 5414 33148 5466
rect 33148 5414 33160 5466
rect 33160 5414 33174 5466
rect 33198 5414 33212 5466
rect 33212 5414 33224 5466
rect 33224 5414 33254 5466
rect 33278 5414 33288 5466
rect 33288 5414 33334 5466
rect 33038 5412 33094 5414
rect 33118 5412 33174 5414
rect 33198 5412 33254 5414
rect 33278 5412 33334 5414
rect 33038 4378 33094 4380
rect 33118 4378 33174 4380
rect 33198 4378 33254 4380
rect 33278 4378 33334 4380
rect 33038 4326 33084 4378
rect 33084 4326 33094 4378
rect 33118 4326 33148 4378
rect 33148 4326 33160 4378
rect 33160 4326 33174 4378
rect 33198 4326 33212 4378
rect 33212 4326 33224 4378
rect 33224 4326 33254 4378
rect 33278 4326 33288 4378
rect 33288 4326 33334 4378
rect 33038 4324 33094 4326
rect 33118 4324 33174 4326
rect 33198 4324 33254 4326
rect 33278 4324 33334 4326
rect 32310 2796 32312 2816
rect 32312 2796 32364 2816
rect 32364 2796 32366 2816
rect 32310 2760 32366 2796
rect 33038 3290 33094 3292
rect 33118 3290 33174 3292
rect 33198 3290 33254 3292
rect 33278 3290 33334 3292
rect 33038 3238 33084 3290
rect 33084 3238 33094 3290
rect 33118 3238 33148 3290
rect 33148 3238 33160 3290
rect 33160 3238 33174 3290
rect 33198 3238 33212 3290
rect 33212 3238 33224 3290
rect 33224 3238 33254 3290
rect 33278 3238 33288 3290
rect 33288 3238 33334 3290
rect 33038 3236 33094 3238
rect 33118 3236 33174 3238
rect 33198 3236 33254 3238
rect 33278 3236 33334 3238
rect 33322 2372 33378 2408
rect 33322 2352 33324 2372
rect 33324 2352 33376 2372
rect 33376 2352 33378 2372
rect 33038 2202 33094 2204
rect 33118 2202 33174 2204
rect 33198 2202 33254 2204
rect 33278 2202 33334 2204
rect 33038 2150 33084 2202
rect 33084 2150 33094 2202
rect 33118 2150 33148 2202
rect 33148 2150 33160 2202
rect 33160 2150 33174 2202
rect 33198 2150 33212 2202
rect 33212 2150 33224 2202
rect 33224 2150 33254 2202
rect 33278 2150 33288 2202
rect 33288 2150 33334 2202
rect 33038 2148 33094 2150
rect 33118 2148 33174 2150
rect 33198 2148 33254 2150
rect 33278 2148 33334 2150
rect 34794 992 34850 1048
rect 43732 7642 43788 7644
rect 43812 7642 43868 7644
rect 43892 7642 43948 7644
rect 43972 7642 44028 7644
rect 43732 7590 43778 7642
rect 43778 7590 43788 7642
rect 43812 7590 43842 7642
rect 43842 7590 43854 7642
rect 43854 7590 43868 7642
rect 43892 7590 43906 7642
rect 43906 7590 43918 7642
rect 43918 7590 43948 7642
rect 43972 7590 43982 7642
rect 43982 7590 44028 7642
rect 43732 7588 43788 7590
rect 43812 7588 43868 7590
rect 43892 7588 43948 7590
rect 43972 7588 44028 7590
rect 38385 7098 38441 7100
rect 38465 7098 38521 7100
rect 38545 7098 38601 7100
rect 38625 7098 38681 7100
rect 38385 7046 38431 7098
rect 38431 7046 38441 7098
rect 38465 7046 38495 7098
rect 38495 7046 38507 7098
rect 38507 7046 38521 7098
rect 38545 7046 38559 7098
rect 38559 7046 38571 7098
rect 38571 7046 38601 7098
rect 38625 7046 38635 7098
rect 38635 7046 38681 7098
rect 38385 7044 38441 7046
rect 38465 7044 38521 7046
rect 38545 7044 38601 7046
rect 38625 7044 38681 7046
rect 36358 2796 36360 2816
rect 36360 2796 36412 2816
rect 36412 2796 36414 2816
rect 36358 2760 36414 2796
rect 38385 6010 38441 6012
rect 38465 6010 38521 6012
rect 38545 6010 38601 6012
rect 38625 6010 38681 6012
rect 38385 5958 38431 6010
rect 38431 5958 38441 6010
rect 38465 5958 38495 6010
rect 38495 5958 38507 6010
rect 38507 5958 38521 6010
rect 38545 5958 38559 6010
rect 38559 5958 38571 6010
rect 38571 5958 38601 6010
rect 38625 5958 38635 6010
rect 38635 5958 38681 6010
rect 38385 5956 38441 5958
rect 38465 5956 38521 5958
rect 38545 5956 38601 5958
rect 38625 5956 38681 5958
rect 37830 2624 37886 2680
rect 38385 4922 38441 4924
rect 38465 4922 38521 4924
rect 38545 4922 38601 4924
rect 38625 4922 38681 4924
rect 38385 4870 38431 4922
rect 38431 4870 38441 4922
rect 38465 4870 38495 4922
rect 38495 4870 38507 4922
rect 38507 4870 38521 4922
rect 38545 4870 38559 4922
rect 38559 4870 38571 4922
rect 38571 4870 38601 4922
rect 38625 4870 38635 4922
rect 38635 4870 38681 4922
rect 38385 4868 38441 4870
rect 38465 4868 38521 4870
rect 38545 4868 38601 4870
rect 38625 4868 38681 4870
rect 38385 3834 38441 3836
rect 38465 3834 38521 3836
rect 38545 3834 38601 3836
rect 38625 3834 38681 3836
rect 38385 3782 38431 3834
rect 38431 3782 38441 3834
rect 38465 3782 38495 3834
rect 38495 3782 38507 3834
rect 38507 3782 38521 3834
rect 38545 3782 38559 3834
rect 38559 3782 38571 3834
rect 38571 3782 38601 3834
rect 38625 3782 38635 3834
rect 38635 3782 38681 3834
rect 38385 3780 38441 3782
rect 38465 3780 38521 3782
rect 38545 3780 38601 3782
rect 38625 3780 38681 3782
rect 38385 2746 38441 2748
rect 38465 2746 38521 2748
rect 38545 2746 38601 2748
rect 38625 2746 38681 2748
rect 38385 2694 38431 2746
rect 38431 2694 38441 2746
rect 38465 2694 38495 2746
rect 38495 2694 38507 2746
rect 38507 2694 38521 2746
rect 38545 2694 38559 2746
rect 38559 2694 38571 2746
rect 38571 2694 38601 2746
rect 38625 2694 38635 2746
rect 38635 2694 38681 2746
rect 38385 2692 38441 2694
rect 38465 2692 38521 2694
rect 38545 2692 38601 2694
rect 38625 2692 38681 2694
rect 43732 6554 43788 6556
rect 43812 6554 43868 6556
rect 43892 6554 43948 6556
rect 43972 6554 44028 6556
rect 43732 6502 43778 6554
rect 43778 6502 43788 6554
rect 43812 6502 43842 6554
rect 43842 6502 43854 6554
rect 43854 6502 43868 6554
rect 43892 6502 43906 6554
rect 43906 6502 43918 6554
rect 43918 6502 43948 6554
rect 43972 6502 43982 6554
rect 43982 6502 44028 6554
rect 43732 6500 43788 6502
rect 43812 6500 43868 6502
rect 43892 6500 43948 6502
rect 43972 6500 44028 6502
rect 43732 5466 43788 5468
rect 43812 5466 43868 5468
rect 43892 5466 43948 5468
rect 43972 5466 44028 5468
rect 43732 5414 43778 5466
rect 43778 5414 43788 5466
rect 43812 5414 43842 5466
rect 43842 5414 43854 5466
rect 43854 5414 43868 5466
rect 43892 5414 43906 5466
rect 43906 5414 43918 5466
rect 43918 5414 43948 5466
rect 43972 5414 43982 5466
rect 43982 5414 44028 5466
rect 43732 5412 43788 5414
rect 43812 5412 43868 5414
rect 43892 5412 43948 5414
rect 43972 5412 44028 5414
rect 43732 4378 43788 4380
rect 43812 4378 43868 4380
rect 43892 4378 43948 4380
rect 43972 4378 44028 4380
rect 43732 4326 43778 4378
rect 43778 4326 43788 4378
rect 43812 4326 43842 4378
rect 43842 4326 43854 4378
rect 43854 4326 43868 4378
rect 43892 4326 43906 4378
rect 43906 4326 43918 4378
rect 43918 4326 43948 4378
rect 43972 4326 43982 4378
rect 43982 4326 44028 4378
rect 43732 4324 43788 4326
rect 43812 4324 43868 4326
rect 43892 4324 43948 4326
rect 43972 4324 44028 4326
rect 43732 3290 43788 3292
rect 43812 3290 43868 3292
rect 43892 3290 43948 3292
rect 43972 3290 44028 3292
rect 43732 3238 43778 3290
rect 43778 3238 43788 3290
rect 43812 3238 43842 3290
rect 43842 3238 43854 3290
rect 43854 3238 43868 3290
rect 43892 3238 43906 3290
rect 43906 3238 43918 3290
rect 43918 3238 43948 3290
rect 43972 3238 43982 3290
rect 43982 3238 44028 3290
rect 43732 3236 43788 3238
rect 43812 3236 43868 3238
rect 43892 3236 43948 3238
rect 43972 3236 44028 3238
rect 43732 2202 43788 2204
rect 43812 2202 43868 2204
rect 43892 2202 43948 2204
rect 43972 2202 44028 2204
rect 43732 2150 43778 2202
rect 43778 2150 43788 2202
rect 43812 2150 43842 2202
rect 43842 2150 43854 2202
rect 43854 2150 43868 2202
rect 43892 2150 43906 2202
rect 43906 2150 43918 2202
rect 43918 2150 43948 2202
rect 43972 2150 43982 2202
rect 43982 2150 44028 2202
rect 43732 2148 43788 2150
rect 43812 2148 43868 2150
rect 43892 2148 43948 2150
rect 43972 2148 44028 2150
<< metal3 >>
rect 11640 7648 11956 7649
rect 11640 7584 11646 7648
rect 11710 7584 11726 7648
rect 11790 7584 11806 7648
rect 11870 7584 11886 7648
rect 11950 7584 11956 7648
rect 11640 7583 11956 7584
rect 22334 7648 22650 7649
rect 22334 7584 22340 7648
rect 22404 7584 22420 7648
rect 22484 7584 22500 7648
rect 22564 7584 22580 7648
rect 22644 7584 22650 7648
rect 22334 7583 22650 7584
rect 33028 7648 33344 7649
rect 33028 7584 33034 7648
rect 33098 7584 33114 7648
rect 33178 7584 33194 7648
rect 33258 7584 33274 7648
rect 33338 7584 33344 7648
rect 33028 7583 33344 7584
rect 43722 7648 44038 7649
rect 43722 7584 43728 7648
rect 43792 7584 43808 7648
rect 43872 7584 43888 7648
rect 43952 7584 43968 7648
rect 44032 7584 44038 7648
rect 43722 7583 44038 7584
rect 6293 7104 6609 7105
rect 6293 7040 6299 7104
rect 6363 7040 6379 7104
rect 6443 7040 6459 7104
rect 6523 7040 6539 7104
rect 6603 7040 6609 7104
rect 6293 7039 6609 7040
rect 16987 7104 17303 7105
rect 16987 7040 16993 7104
rect 17057 7040 17073 7104
rect 17137 7040 17153 7104
rect 17217 7040 17233 7104
rect 17297 7040 17303 7104
rect 16987 7039 17303 7040
rect 27681 7104 27997 7105
rect 27681 7040 27687 7104
rect 27751 7040 27767 7104
rect 27831 7040 27847 7104
rect 27911 7040 27927 7104
rect 27991 7040 27997 7104
rect 27681 7039 27997 7040
rect 38375 7104 38691 7105
rect 38375 7040 38381 7104
rect 38445 7040 38461 7104
rect 38525 7040 38541 7104
rect 38605 7040 38621 7104
rect 38685 7040 38691 7104
rect 38375 7039 38691 7040
rect 11640 6560 11956 6561
rect 11640 6496 11646 6560
rect 11710 6496 11726 6560
rect 11790 6496 11806 6560
rect 11870 6496 11886 6560
rect 11950 6496 11956 6560
rect 11640 6495 11956 6496
rect 22334 6560 22650 6561
rect 22334 6496 22340 6560
rect 22404 6496 22420 6560
rect 22484 6496 22500 6560
rect 22564 6496 22580 6560
rect 22644 6496 22650 6560
rect 22334 6495 22650 6496
rect 33028 6560 33344 6561
rect 33028 6496 33034 6560
rect 33098 6496 33114 6560
rect 33178 6496 33194 6560
rect 33258 6496 33274 6560
rect 33338 6496 33344 6560
rect 33028 6495 33344 6496
rect 43722 6560 44038 6561
rect 43722 6496 43728 6560
rect 43792 6496 43808 6560
rect 43872 6496 43888 6560
rect 43952 6496 43968 6560
rect 44032 6496 44038 6560
rect 43722 6495 44038 6496
rect 6293 6016 6609 6017
rect 6293 5952 6299 6016
rect 6363 5952 6379 6016
rect 6443 5952 6459 6016
rect 6523 5952 6539 6016
rect 6603 5952 6609 6016
rect 6293 5951 6609 5952
rect 16987 6016 17303 6017
rect 16987 5952 16993 6016
rect 17057 5952 17073 6016
rect 17137 5952 17153 6016
rect 17217 5952 17233 6016
rect 17297 5952 17303 6016
rect 16987 5951 17303 5952
rect 27681 6016 27997 6017
rect 27681 5952 27687 6016
rect 27751 5952 27767 6016
rect 27831 5952 27847 6016
rect 27911 5952 27927 6016
rect 27991 5952 27997 6016
rect 27681 5951 27997 5952
rect 38375 6016 38691 6017
rect 38375 5952 38381 6016
rect 38445 5952 38461 6016
rect 38525 5952 38541 6016
rect 38605 5952 38621 6016
rect 38685 5952 38691 6016
rect 38375 5951 38691 5952
rect 16481 5674 16547 5677
rect 36854 5674 36860 5676
rect 16481 5672 36860 5674
rect 16481 5616 16486 5672
rect 16542 5616 36860 5672
rect 16481 5614 36860 5616
rect 16481 5611 16547 5614
rect 36854 5612 36860 5614
rect 36924 5612 36930 5676
rect 11640 5472 11956 5473
rect 11640 5408 11646 5472
rect 11710 5408 11726 5472
rect 11790 5408 11806 5472
rect 11870 5408 11886 5472
rect 11950 5408 11956 5472
rect 11640 5407 11956 5408
rect 22334 5472 22650 5473
rect 22334 5408 22340 5472
rect 22404 5408 22420 5472
rect 22484 5408 22500 5472
rect 22564 5408 22580 5472
rect 22644 5408 22650 5472
rect 22334 5407 22650 5408
rect 33028 5472 33344 5473
rect 33028 5408 33034 5472
rect 33098 5408 33114 5472
rect 33178 5408 33194 5472
rect 33258 5408 33274 5472
rect 33338 5408 33344 5472
rect 33028 5407 33344 5408
rect 43722 5472 44038 5473
rect 43722 5408 43728 5472
rect 43792 5408 43808 5472
rect 43872 5408 43888 5472
rect 43952 5408 43968 5472
rect 44032 5408 44038 5472
rect 43722 5407 44038 5408
rect 6293 4928 6609 4929
rect 6293 4864 6299 4928
rect 6363 4864 6379 4928
rect 6443 4864 6459 4928
rect 6523 4864 6539 4928
rect 6603 4864 6609 4928
rect 6293 4863 6609 4864
rect 16987 4928 17303 4929
rect 16987 4864 16993 4928
rect 17057 4864 17073 4928
rect 17137 4864 17153 4928
rect 17217 4864 17233 4928
rect 17297 4864 17303 4928
rect 16987 4863 17303 4864
rect 27681 4928 27997 4929
rect 27681 4864 27687 4928
rect 27751 4864 27767 4928
rect 27831 4864 27847 4928
rect 27911 4864 27927 4928
rect 27991 4864 27997 4928
rect 27681 4863 27997 4864
rect 38375 4928 38691 4929
rect 38375 4864 38381 4928
rect 38445 4864 38461 4928
rect 38525 4864 38541 4928
rect 38605 4864 38621 4928
rect 38685 4864 38691 4928
rect 38375 4863 38691 4864
rect 7925 4722 7991 4725
rect 22093 4722 22159 4725
rect 7925 4720 22159 4722
rect 7925 4664 7930 4720
rect 7986 4664 22098 4720
rect 22154 4664 22159 4720
rect 7925 4662 22159 4664
rect 7925 4659 7991 4662
rect 22093 4659 22159 4662
rect 8201 4586 8267 4589
rect 22001 4586 22067 4589
rect 8201 4584 22067 4586
rect 8201 4528 8206 4584
rect 8262 4528 22006 4584
rect 22062 4528 22067 4584
rect 8201 4526 22067 4528
rect 8201 4523 8267 4526
rect 22001 4523 22067 4526
rect 11640 4384 11956 4385
rect 11640 4320 11646 4384
rect 11710 4320 11726 4384
rect 11790 4320 11806 4384
rect 11870 4320 11886 4384
rect 11950 4320 11956 4384
rect 11640 4319 11956 4320
rect 22334 4384 22650 4385
rect 22334 4320 22340 4384
rect 22404 4320 22420 4384
rect 22484 4320 22500 4384
rect 22564 4320 22580 4384
rect 22644 4320 22650 4384
rect 22334 4319 22650 4320
rect 33028 4384 33344 4385
rect 33028 4320 33034 4384
rect 33098 4320 33114 4384
rect 33178 4320 33194 4384
rect 33258 4320 33274 4384
rect 33338 4320 33344 4384
rect 33028 4319 33344 4320
rect 43722 4384 44038 4385
rect 43722 4320 43728 4384
rect 43792 4320 43808 4384
rect 43872 4320 43888 4384
rect 43952 4320 43968 4384
rect 44032 4320 44038 4384
rect 43722 4319 44038 4320
rect 11973 4042 12039 4045
rect 24945 4042 25011 4045
rect 11973 4040 25011 4042
rect 11973 3984 11978 4040
rect 12034 3984 24950 4040
rect 25006 3984 25011 4040
rect 11973 3982 25011 3984
rect 11973 3979 12039 3982
rect 24945 3979 25011 3982
rect 6293 3840 6609 3841
rect 6293 3776 6299 3840
rect 6363 3776 6379 3840
rect 6443 3776 6459 3840
rect 6523 3776 6539 3840
rect 6603 3776 6609 3840
rect 6293 3775 6609 3776
rect 16987 3840 17303 3841
rect 16987 3776 16993 3840
rect 17057 3776 17073 3840
rect 17137 3776 17153 3840
rect 17217 3776 17233 3840
rect 17297 3776 17303 3840
rect 16987 3775 17303 3776
rect 27681 3840 27997 3841
rect 27681 3776 27687 3840
rect 27751 3776 27767 3840
rect 27831 3776 27847 3840
rect 27911 3776 27927 3840
rect 27991 3776 27997 3840
rect 27681 3775 27997 3776
rect 38375 3840 38691 3841
rect 38375 3776 38381 3840
rect 38445 3776 38461 3840
rect 38525 3776 38541 3840
rect 38605 3776 38621 3840
rect 38685 3776 38691 3840
rect 38375 3775 38691 3776
rect 19149 3770 19215 3773
rect 26233 3770 26299 3773
rect 19149 3768 26299 3770
rect 19149 3712 19154 3768
rect 19210 3712 26238 3768
rect 26294 3712 26299 3768
rect 19149 3710 26299 3712
rect 19149 3707 19215 3710
rect 26233 3707 26299 3710
rect 11053 3634 11119 3637
rect 27613 3634 27679 3637
rect 11053 3632 27679 3634
rect 11053 3576 11058 3632
rect 11114 3576 27618 3632
rect 27674 3576 27679 3632
rect 11053 3574 27679 3576
rect 11053 3571 11119 3574
rect 27613 3571 27679 3574
rect 12525 3498 12591 3501
rect 26509 3498 26575 3501
rect 12525 3496 26575 3498
rect 12525 3440 12530 3496
rect 12586 3440 26514 3496
rect 26570 3440 26575 3496
rect 12525 3438 26575 3440
rect 12525 3435 12591 3438
rect 26509 3435 26575 3438
rect 11640 3296 11956 3297
rect 11640 3232 11646 3296
rect 11710 3232 11726 3296
rect 11790 3232 11806 3296
rect 11870 3232 11886 3296
rect 11950 3232 11956 3296
rect 11640 3231 11956 3232
rect 22334 3296 22650 3297
rect 22334 3232 22340 3296
rect 22404 3232 22420 3296
rect 22484 3232 22500 3296
rect 22564 3232 22580 3296
rect 22644 3232 22650 3296
rect 22334 3231 22650 3232
rect 33028 3296 33344 3297
rect 33028 3232 33034 3296
rect 33098 3232 33114 3296
rect 33178 3232 33194 3296
rect 33258 3232 33274 3296
rect 33338 3232 33344 3296
rect 33028 3231 33344 3232
rect 43722 3296 44038 3297
rect 43722 3232 43728 3296
rect 43792 3232 43808 3296
rect 43872 3232 43888 3296
rect 43952 3232 43968 3296
rect 44032 3232 44038 3296
rect 43722 3231 44038 3232
rect 18229 3226 18295 3229
rect 18229 3224 22110 3226
rect 18229 3168 18234 3224
rect 18290 3168 22110 3224
rect 18229 3166 22110 3168
rect 18229 3163 18295 3166
rect 8753 3090 8819 3093
rect 21357 3090 21423 3093
rect 8753 3088 21423 3090
rect 8753 3032 8758 3088
rect 8814 3032 21362 3088
rect 21418 3032 21423 3088
rect 8753 3030 21423 3032
rect 22050 3090 22110 3166
rect 28993 3090 29059 3093
rect 22050 3088 29059 3090
rect 22050 3032 28998 3088
rect 29054 3032 29059 3088
rect 22050 3030 29059 3032
rect 8753 3027 8819 3030
rect 21357 3027 21423 3030
rect 28993 3027 29059 3030
rect 18321 2954 18387 2957
rect 29085 2954 29151 2957
rect 18321 2952 29151 2954
rect 18321 2896 18326 2952
rect 18382 2896 29090 2952
rect 29146 2896 29151 2952
rect 18321 2894 29151 2896
rect 18321 2891 18387 2894
rect 29085 2891 29151 2894
rect 26785 2818 26851 2821
rect 20670 2816 26851 2818
rect 20670 2760 26790 2816
rect 26846 2760 26851 2816
rect 20670 2758 26851 2760
rect 6293 2752 6609 2753
rect 6293 2688 6299 2752
rect 6363 2688 6379 2752
rect 6443 2688 6459 2752
rect 6523 2688 6539 2752
rect 6603 2688 6609 2752
rect 6293 2687 6609 2688
rect 16987 2752 17303 2753
rect 16987 2688 16993 2752
rect 17057 2688 17073 2752
rect 17137 2688 17153 2752
rect 17217 2688 17233 2752
rect 17297 2688 17303 2752
rect 16987 2687 17303 2688
rect 20670 2682 20730 2758
rect 26785 2755 26851 2758
rect 30230 2756 30236 2820
rect 30300 2818 30306 2820
rect 32305 2818 32371 2821
rect 30300 2816 32371 2818
rect 30300 2760 32310 2816
rect 32366 2760 32371 2816
rect 30300 2758 32371 2760
rect 30300 2756 30306 2758
rect 32305 2755 32371 2758
rect 36118 2756 36124 2820
rect 36188 2818 36194 2820
rect 36353 2818 36419 2821
rect 36188 2816 36419 2818
rect 36188 2760 36358 2816
rect 36414 2760 36419 2816
rect 36188 2758 36419 2760
rect 36188 2756 36194 2758
rect 36353 2755 36419 2758
rect 27681 2752 27997 2753
rect 27681 2688 27687 2752
rect 27751 2688 27767 2752
rect 27831 2688 27847 2752
rect 27911 2688 27927 2752
rect 27991 2688 27997 2752
rect 27681 2687 27997 2688
rect 38375 2752 38691 2753
rect 38375 2688 38381 2752
rect 38445 2688 38461 2752
rect 38525 2688 38541 2752
rect 38605 2688 38621 2752
rect 38685 2688 38691 2752
rect 38375 2687 38691 2688
rect 18646 2622 20730 2682
rect 18229 2410 18295 2413
rect 11102 2408 18295 2410
rect 11102 2352 18234 2408
rect 18290 2352 18295 2408
rect 11102 2350 18295 2352
rect 11102 2277 11162 2350
rect 18229 2347 18295 2350
rect 11053 2272 11162 2277
rect 11053 2216 11058 2272
rect 11114 2216 11162 2272
rect 11053 2214 11162 2216
rect 12249 2274 12315 2277
rect 18646 2274 18706 2622
rect 36854 2620 36860 2684
rect 36924 2682 36930 2684
rect 37825 2682 37891 2685
rect 36924 2680 37891 2682
rect 36924 2624 37830 2680
rect 37886 2624 37891 2680
rect 36924 2622 37891 2624
rect 36924 2620 36930 2622
rect 37825 2619 37891 2622
rect 18873 2546 18939 2549
rect 27889 2546 27955 2549
rect 18873 2544 27955 2546
rect 18873 2488 18878 2544
rect 18934 2488 27894 2544
rect 27950 2488 27955 2544
rect 18873 2486 27955 2488
rect 18873 2483 18939 2486
rect 27889 2483 27955 2486
rect 33317 2410 33383 2413
rect 12249 2272 18706 2274
rect 12249 2216 12254 2272
rect 12310 2216 18706 2272
rect 12249 2214 18706 2216
rect 22050 2408 33383 2410
rect 22050 2352 33322 2408
rect 33378 2352 33383 2408
rect 22050 2350 33383 2352
rect 11053 2211 11119 2214
rect 12249 2211 12315 2214
rect 11640 2208 11956 2209
rect 11640 2144 11646 2208
rect 11710 2144 11726 2208
rect 11790 2144 11806 2208
rect 11870 2144 11886 2208
rect 11950 2144 11956 2208
rect 11640 2143 11956 2144
rect 12157 2138 12223 2141
rect 18321 2138 18387 2141
rect 12157 2136 18387 2138
rect 12157 2080 12162 2136
rect 12218 2080 18326 2136
rect 18382 2080 18387 2136
rect 12157 2078 18387 2080
rect 12157 2075 12223 2078
rect 18321 2075 18387 2078
rect 19149 2002 19215 2005
rect 22050 2002 22110 2350
rect 33317 2347 33383 2350
rect 22334 2208 22650 2209
rect 22334 2144 22340 2208
rect 22404 2144 22420 2208
rect 22484 2144 22500 2208
rect 22564 2144 22580 2208
rect 22644 2144 22650 2208
rect 22334 2143 22650 2144
rect 33028 2208 33344 2209
rect 33028 2144 33034 2208
rect 33098 2144 33114 2208
rect 33178 2144 33194 2208
rect 33258 2144 33274 2208
rect 33338 2144 33344 2208
rect 33028 2143 33344 2144
rect 43722 2208 44038 2209
rect 43722 2144 43728 2208
rect 43792 2144 43808 2208
rect 43872 2144 43888 2208
rect 43952 2144 43968 2208
rect 44032 2144 44038 2208
rect 43722 2143 44038 2144
rect 27153 2002 27219 2005
rect 19149 2000 22110 2002
rect 19149 1944 19154 2000
rect 19210 1944 22110 2000
rect 19149 1942 22110 1944
rect 24534 2000 27219 2002
rect 24534 1944 27158 2000
rect 27214 1944 27219 2000
rect 24534 1942 27219 1944
rect 19149 1939 19215 1942
rect 13261 1866 13327 1869
rect 24534 1866 24594 1942
rect 27153 1939 27219 1942
rect 13261 1864 24594 1866
rect 13261 1808 13266 1864
rect 13322 1808 24594 1864
rect 13261 1806 24594 1808
rect 13261 1803 13327 1806
rect 17309 1730 17375 1733
rect 30373 1730 30439 1733
rect 17309 1728 30439 1730
rect 17309 1672 17314 1728
rect 17370 1672 30378 1728
rect 30434 1672 30439 1728
rect 17309 1670 30439 1672
rect 17309 1667 17375 1670
rect 30373 1667 30439 1670
rect 10501 1594 10567 1597
rect 28533 1594 28599 1597
rect 10501 1592 28599 1594
rect 10501 1536 10506 1592
rect 10562 1536 28538 1592
rect 28594 1536 28599 1592
rect 10501 1534 28599 1536
rect 10501 1531 10567 1534
rect 28533 1531 28599 1534
rect 9397 1458 9463 1461
rect 21081 1458 21147 1461
rect 9397 1456 21147 1458
rect 9397 1400 9402 1456
rect 9458 1400 21086 1456
rect 21142 1400 21147 1456
rect 9397 1398 21147 1400
rect 9397 1395 9463 1398
rect 21081 1395 21147 1398
rect 19149 1322 19215 1325
rect 30230 1322 30236 1324
rect 19149 1320 30236 1322
rect 19149 1264 19154 1320
rect 19210 1264 30236 1320
rect 19149 1262 30236 1264
rect 19149 1259 19215 1262
rect 30230 1260 30236 1262
rect 30300 1260 30306 1324
rect 10777 1186 10843 1189
rect 28441 1186 28507 1189
rect 10777 1184 28507 1186
rect 10777 1128 10782 1184
rect 10838 1128 28446 1184
rect 28502 1128 28507 1184
rect 10777 1126 28507 1128
rect 10777 1123 10843 1126
rect 28441 1123 28507 1126
rect 16665 1050 16731 1053
rect 34789 1050 34855 1053
rect 16665 1048 34855 1050
rect 16665 992 16670 1048
rect 16726 992 34794 1048
rect 34850 992 34855 1048
rect 16665 990 34855 992
rect 16665 987 16731 990
rect 34789 987 34855 990
rect 14825 914 14891 917
rect 36118 914 36124 916
rect 14825 912 36124 914
rect 14825 856 14830 912
rect 14886 856 36124 912
rect 14825 854 36124 856
rect 14825 851 14891 854
rect 36118 852 36124 854
rect 36188 852 36194 916
<< via3 >>
rect 11646 7644 11710 7648
rect 11646 7588 11650 7644
rect 11650 7588 11706 7644
rect 11706 7588 11710 7644
rect 11646 7584 11710 7588
rect 11726 7644 11790 7648
rect 11726 7588 11730 7644
rect 11730 7588 11786 7644
rect 11786 7588 11790 7644
rect 11726 7584 11790 7588
rect 11806 7644 11870 7648
rect 11806 7588 11810 7644
rect 11810 7588 11866 7644
rect 11866 7588 11870 7644
rect 11806 7584 11870 7588
rect 11886 7644 11950 7648
rect 11886 7588 11890 7644
rect 11890 7588 11946 7644
rect 11946 7588 11950 7644
rect 11886 7584 11950 7588
rect 22340 7644 22404 7648
rect 22340 7588 22344 7644
rect 22344 7588 22400 7644
rect 22400 7588 22404 7644
rect 22340 7584 22404 7588
rect 22420 7644 22484 7648
rect 22420 7588 22424 7644
rect 22424 7588 22480 7644
rect 22480 7588 22484 7644
rect 22420 7584 22484 7588
rect 22500 7644 22564 7648
rect 22500 7588 22504 7644
rect 22504 7588 22560 7644
rect 22560 7588 22564 7644
rect 22500 7584 22564 7588
rect 22580 7644 22644 7648
rect 22580 7588 22584 7644
rect 22584 7588 22640 7644
rect 22640 7588 22644 7644
rect 22580 7584 22644 7588
rect 33034 7644 33098 7648
rect 33034 7588 33038 7644
rect 33038 7588 33094 7644
rect 33094 7588 33098 7644
rect 33034 7584 33098 7588
rect 33114 7644 33178 7648
rect 33114 7588 33118 7644
rect 33118 7588 33174 7644
rect 33174 7588 33178 7644
rect 33114 7584 33178 7588
rect 33194 7644 33258 7648
rect 33194 7588 33198 7644
rect 33198 7588 33254 7644
rect 33254 7588 33258 7644
rect 33194 7584 33258 7588
rect 33274 7644 33338 7648
rect 33274 7588 33278 7644
rect 33278 7588 33334 7644
rect 33334 7588 33338 7644
rect 33274 7584 33338 7588
rect 43728 7644 43792 7648
rect 43728 7588 43732 7644
rect 43732 7588 43788 7644
rect 43788 7588 43792 7644
rect 43728 7584 43792 7588
rect 43808 7644 43872 7648
rect 43808 7588 43812 7644
rect 43812 7588 43868 7644
rect 43868 7588 43872 7644
rect 43808 7584 43872 7588
rect 43888 7644 43952 7648
rect 43888 7588 43892 7644
rect 43892 7588 43948 7644
rect 43948 7588 43952 7644
rect 43888 7584 43952 7588
rect 43968 7644 44032 7648
rect 43968 7588 43972 7644
rect 43972 7588 44028 7644
rect 44028 7588 44032 7644
rect 43968 7584 44032 7588
rect 6299 7100 6363 7104
rect 6299 7044 6303 7100
rect 6303 7044 6359 7100
rect 6359 7044 6363 7100
rect 6299 7040 6363 7044
rect 6379 7100 6443 7104
rect 6379 7044 6383 7100
rect 6383 7044 6439 7100
rect 6439 7044 6443 7100
rect 6379 7040 6443 7044
rect 6459 7100 6523 7104
rect 6459 7044 6463 7100
rect 6463 7044 6519 7100
rect 6519 7044 6523 7100
rect 6459 7040 6523 7044
rect 6539 7100 6603 7104
rect 6539 7044 6543 7100
rect 6543 7044 6599 7100
rect 6599 7044 6603 7100
rect 6539 7040 6603 7044
rect 16993 7100 17057 7104
rect 16993 7044 16997 7100
rect 16997 7044 17053 7100
rect 17053 7044 17057 7100
rect 16993 7040 17057 7044
rect 17073 7100 17137 7104
rect 17073 7044 17077 7100
rect 17077 7044 17133 7100
rect 17133 7044 17137 7100
rect 17073 7040 17137 7044
rect 17153 7100 17217 7104
rect 17153 7044 17157 7100
rect 17157 7044 17213 7100
rect 17213 7044 17217 7100
rect 17153 7040 17217 7044
rect 17233 7100 17297 7104
rect 17233 7044 17237 7100
rect 17237 7044 17293 7100
rect 17293 7044 17297 7100
rect 17233 7040 17297 7044
rect 27687 7100 27751 7104
rect 27687 7044 27691 7100
rect 27691 7044 27747 7100
rect 27747 7044 27751 7100
rect 27687 7040 27751 7044
rect 27767 7100 27831 7104
rect 27767 7044 27771 7100
rect 27771 7044 27827 7100
rect 27827 7044 27831 7100
rect 27767 7040 27831 7044
rect 27847 7100 27911 7104
rect 27847 7044 27851 7100
rect 27851 7044 27907 7100
rect 27907 7044 27911 7100
rect 27847 7040 27911 7044
rect 27927 7100 27991 7104
rect 27927 7044 27931 7100
rect 27931 7044 27987 7100
rect 27987 7044 27991 7100
rect 27927 7040 27991 7044
rect 38381 7100 38445 7104
rect 38381 7044 38385 7100
rect 38385 7044 38441 7100
rect 38441 7044 38445 7100
rect 38381 7040 38445 7044
rect 38461 7100 38525 7104
rect 38461 7044 38465 7100
rect 38465 7044 38521 7100
rect 38521 7044 38525 7100
rect 38461 7040 38525 7044
rect 38541 7100 38605 7104
rect 38541 7044 38545 7100
rect 38545 7044 38601 7100
rect 38601 7044 38605 7100
rect 38541 7040 38605 7044
rect 38621 7100 38685 7104
rect 38621 7044 38625 7100
rect 38625 7044 38681 7100
rect 38681 7044 38685 7100
rect 38621 7040 38685 7044
rect 11646 6556 11710 6560
rect 11646 6500 11650 6556
rect 11650 6500 11706 6556
rect 11706 6500 11710 6556
rect 11646 6496 11710 6500
rect 11726 6556 11790 6560
rect 11726 6500 11730 6556
rect 11730 6500 11786 6556
rect 11786 6500 11790 6556
rect 11726 6496 11790 6500
rect 11806 6556 11870 6560
rect 11806 6500 11810 6556
rect 11810 6500 11866 6556
rect 11866 6500 11870 6556
rect 11806 6496 11870 6500
rect 11886 6556 11950 6560
rect 11886 6500 11890 6556
rect 11890 6500 11946 6556
rect 11946 6500 11950 6556
rect 11886 6496 11950 6500
rect 22340 6556 22404 6560
rect 22340 6500 22344 6556
rect 22344 6500 22400 6556
rect 22400 6500 22404 6556
rect 22340 6496 22404 6500
rect 22420 6556 22484 6560
rect 22420 6500 22424 6556
rect 22424 6500 22480 6556
rect 22480 6500 22484 6556
rect 22420 6496 22484 6500
rect 22500 6556 22564 6560
rect 22500 6500 22504 6556
rect 22504 6500 22560 6556
rect 22560 6500 22564 6556
rect 22500 6496 22564 6500
rect 22580 6556 22644 6560
rect 22580 6500 22584 6556
rect 22584 6500 22640 6556
rect 22640 6500 22644 6556
rect 22580 6496 22644 6500
rect 33034 6556 33098 6560
rect 33034 6500 33038 6556
rect 33038 6500 33094 6556
rect 33094 6500 33098 6556
rect 33034 6496 33098 6500
rect 33114 6556 33178 6560
rect 33114 6500 33118 6556
rect 33118 6500 33174 6556
rect 33174 6500 33178 6556
rect 33114 6496 33178 6500
rect 33194 6556 33258 6560
rect 33194 6500 33198 6556
rect 33198 6500 33254 6556
rect 33254 6500 33258 6556
rect 33194 6496 33258 6500
rect 33274 6556 33338 6560
rect 33274 6500 33278 6556
rect 33278 6500 33334 6556
rect 33334 6500 33338 6556
rect 33274 6496 33338 6500
rect 43728 6556 43792 6560
rect 43728 6500 43732 6556
rect 43732 6500 43788 6556
rect 43788 6500 43792 6556
rect 43728 6496 43792 6500
rect 43808 6556 43872 6560
rect 43808 6500 43812 6556
rect 43812 6500 43868 6556
rect 43868 6500 43872 6556
rect 43808 6496 43872 6500
rect 43888 6556 43952 6560
rect 43888 6500 43892 6556
rect 43892 6500 43948 6556
rect 43948 6500 43952 6556
rect 43888 6496 43952 6500
rect 43968 6556 44032 6560
rect 43968 6500 43972 6556
rect 43972 6500 44028 6556
rect 44028 6500 44032 6556
rect 43968 6496 44032 6500
rect 6299 6012 6363 6016
rect 6299 5956 6303 6012
rect 6303 5956 6359 6012
rect 6359 5956 6363 6012
rect 6299 5952 6363 5956
rect 6379 6012 6443 6016
rect 6379 5956 6383 6012
rect 6383 5956 6439 6012
rect 6439 5956 6443 6012
rect 6379 5952 6443 5956
rect 6459 6012 6523 6016
rect 6459 5956 6463 6012
rect 6463 5956 6519 6012
rect 6519 5956 6523 6012
rect 6459 5952 6523 5956
rect 6539 6012 6603 6016
rect 6539 5956 6543 6012
rect 6543 5956 6599 6012
rect 6599 5956 6603 6012
rect 6539 5952 6603 5956
rect 16993 6012 17057 6016
rect 16993 5956 16997 6012
rect 16997 5956 17053 6012
rect 17053 5956 17057 6012
rect 16993 5952 17057 5956
rect 17073 6012 17137 6016
rect 17073 5956 17077 6012
rect 17077 5956 17133 6012
rect 17133 5956 17137 6012
rect 17073 5952 17137 5956
rect 17153 6012 17217 6016
rect 17153 5956 17157 6012
rect 17157 5956 17213 6012
rect 17213 5956 17217 6012
rect 17153 5952 17217 5956
rect 17233 6012 17297 6016
rect 17233 5956 17237 6012
rect 17237 5956 17293 6012
rect 17293 5956 17297 6012
rect 17233 5952 17297 5956
rect 27687 6012 27751 6016
rect 27687 5956 27691 6012
rect 27691 5956 27747 6012
rect 27747 5956 27751 6012
rect 27687 5952 27751 5956
rect 27767 6012 27831 6016
rect 27767 5956 27771 6012
rect 27771 5956 27827 6012
rect 27827 5956 27831 6012
rect 27767 5952 27831 5956
rect 27847 6012 27911 6016
rect 27847 5956 27851 6012
rect 27851 5956 27907 6012
rect 27907 5956 27911 6012
rect 27847 5952 27911 5956
rect 27927 6012 27991 6016
rect 27927 5956 27931 6012
rect 27931 5956 27987 6012
rect 27987 5956 27991 6012
rect 27927 5952 27991 5956
rect 38381 6012 38445 6016
rect 38381 5956 38385 6012
rect 38385 5956 38441 6012
rect 38441 5956 38445 6012
rect 38381 5952 38445 5956
rect 38461 6012 38525 6016
rect 38461 5956 38465 6012
rect 38465 5956 38521 6012
rect 38521 5956 38525 6012
rect 38461 5952 38525 5956
rect 38541 6012 38605 6016
rect 38541 5956 38545 6012
rect 38545 5956 38601 6012
rect 38601 5956 38605 6012
rect 38541 5952 38605 5956
rect 38621 6012 38685 6016
rect 38621 5956 38625 6012
rect 38625 5956 38681 6012
rect 38681 5956 38685 6012
rect 38621 5952 38685 5956
rect 36860 5612 36924 5676
rect 11646 5468 11710 5472
rect 11646 5412 11650 5468
rect 11650 5412 11706 5468
rect 11706 5412 11710 5468
rect 11646 5408 11710 5412
rect 11726 5468 11790 5472
rect 11726 5412 11730 5468
rect 11730 5412 11786 5468
rect 11786 5412 11790 5468
rect 11726 5408 11790 5412
rect 11806 5468 11870 5472
rect 11806 5412 11810 5468
rect 11810 5412 11866 5468
rect 11866 5412 11870 5468
rect 11806 5408 11870 5412
rect 11886 5468 11950 5472
rect 11886 5412 11890 5468
rect 11890 5412 11946 5468
rect 11946 5412 11950 5468
rect 11886 5408 11950 5412
rect 22340 5468 22404 5472
rect 22340 5412 22344 5468
rect 22344 5412 22400 5468
rect 22400 5412 22404 5468
rect 22340 5408 22404 5412
rect 22420 5468 22484 5472
rect 22420 5412 22424 5468
rect 22424 5412 22480 5468
rect 22480 5412 22484 5468
rect 22420 5408 22484 5412
rect 22500 5468 22564 5472
rect 22500 5412 22504 5468
rect 22504 5412 22560 5468
rect 22560 5412 22564 5468
rect 22500 5408 22564 5412
rect 22580 5468 22644 5472
rect 22580 5412 22584 5468
rect 22584 5412 22640 5468
rect 22640 5412 22644 5468
rect 22580 5408 22644 5412
rect 33034 5468 33098 5472
rect 33034 5412 33038 5468
rect 33038 5412 33094 5468
rect 33094 5412 33098 5468
rect 33034 5408 33098 5412
rect 33114 5468 33178 5472
rect 33114 5412 33118 5468
rect 33118 5412 33174 5468
rect 33174 5412 33178 5468
rect 33114 5408 33178 5412
rect 33194 5468 33258 5472
rect 33194 5412 33198 5468
rect 33198 5412 33254 5468
rect 33254 5412 33258 5468
rect 33194 5408 33258 5412
rect 33274 5468 33338 5472
rect 33274 5412 33278 5468
rect 33278 5412 33334 5468
rect 33334 5412 33338 5468
rect 33274 5408 33338 5412
rect 43728 5468 43792 5472
rect 43728 5412 43732 5468
rect 43732 5412 43788 5468
rect 43788 5412 43792 5468
rect 43728 5408 43792 5412
rect 43808 5468 43872 5472
rect 43808 5412 43812 5468
rect 43812 5412 43868 5468
rect 43868 5412 43872 5468
rect 43808 5408 43872 5412
rect 43888 5468 43952 5472
rect 43888 5412 43892 5468
rect 43892 5412 43948 5468
rect 43948 5412 43952 5468
rect 43888 5408 43952 5412
rect 43968 5468 44032 5472
rect 43968 5412 43972 5468
rect 43972 5412 44028 5468
rect 44028 5412 44032 5468
rect 43968 5408 44032 5412
rect 6299 4924 6363 4928
rect 6299 4868 6303 4924
rect 6303 4868 6359 4924
rect 6359 4868 6363 4924
rect 6299 4864 6363 4868
rect 6379 4924 6443 4928
rect 6379 4868 6383 4924
rect 6383 4868 6439 4924
rect 6439 4868 6443 4924
rect 6379 4864 6443 4868
rect 6459 4924 6523 4928
rect 6459 4868 6463 4924
rect 6463 4868 6519 4924
rect 6519 4868 6523 4924
rect 6459 4864 6523 4868
rect 6539 4924 6603 4928
rect 6539 4868 6543 4924
rect 6543 4868 6599 4924
rect 6599 4868 6603 4924
rect 6539 4864 6603 4868
rect 16993 4924 17057 4928
rect 16993 4868 16997 4924
rect 16997 4868 17053 4924
rect 17053 4868 17057 4924
rect 16993 4864 17057 4868
rect 17073 4924 17137 4928
rect 17073 4868 17077 4924
rect 17077 4868 17133 4924
rect 17133 4868 17137 4924
rect 17073 4864 17137 4868
rect 17153 4924 17217 4928
rect 17153 4868 17157 4924
rect 17157 4868 17213 4924
rect 17213 4868 17217 4924
rect 17153 4864 17217 4868
rect 17233 4924 17297 4928
rect 17233 4868 17237 4924
rect 17237 4868 17293 4924
rect 17293 4868 17297 4924
rect 17233 4864 17297 4868
rect 27687 4924 27751 4928
rect 27687 4868 27691 4924
rect 27691 4868 27747 4924
rect 27747 4868 27751 4924
rect 27687 4864 27751 4868
rect 27767 4924 27831 4928
rect 27767 4868 27771 4924
rect 27771 4868 27827 4924
rect 27827 4868 27831 4924
rect 27767 4864 27831 4868
rect 27847 4924 27911 4928
rect 27847 4868 27851 4924
rect 27851 4868 27907 4924
rect 27907 4868 27911 4924
rect 27847 4864 27911 4868
rect 27927 4924 27991 4928
rect 27927 4868 27931 4924
rect 27931 4868 27987 4924
rect 27987 4868 27991 4924
rect 27927 4864 27991 4868
rect 38381 4924 38445 4928
rect 38381 4868 38385 4924
rect 38385 4868 38441 4924
rect 38441 4868 38445 4924
rect 38381 4864 38445 4868
rect 38461 4924 38525 4928
rect 38461 4868 38465 4924
rect 38465 4868 38521 4924
rect 38521 4868 38525 4924
rect 38461 4864 38525 4868
rect 38541 4924 38605 4928
rect 38541 4868 38545 4924
rect 38545 4868 38601 4924
rect 38601 4868 38605 4924
rect 38541 4864 38605 4868
rect 38621 4924 38685 4928
rect 38621 4868 38625 4924
rect 38625 4868 38681 4924
rect 38681 4868 38685 4924
rect 38621 4864 38685 4868
rect 11646 4380 11710 4384
rect 11646 4324 11650 4380
rect 11650 4324 11706 4380
rect 11706 4324 11710 4380
rect 11646 4320 11710 4324
rect 11726 4380 11790 4384
rect 11726 4324 11730 4380
rect 11730 4324 11786 4380
rect 11786 4324 11790 4380
rect 11726 4320 11790 4324
rect 11806 4380 11870 4384
rect 11806 4324 11810 4380
rect 11810 4324 11866 4380
rect 11866 4324 11870 4380
rect 11806 4320 11870 4324
rect 11886 4380 11950 4384
rect 11886 4324 11890 4380
rect 11890 4324 11946 4380
rect 11946 4324 11950 4380
rect 11886 4320 11950 4324
rect 22340 4380 22404 4384
rect 22340 4324 22344 4380
rect 22344 4324 22400 4380
rect 22400 4324 22404 4380
rect 22340 4320 22404 4324
rect 22420 4380 22484 4384
rect 22420 4324 22424 4380
rect 22424 4324 22480 4380
rect 22480 4324 22484 4380
rect 22420 4320 22484 4324
rect 22500 4380 22564 4384
rect 22500 4324 22504 4380
rect 22504 4324 22560 4380
rect 22560 4324 22564 4380
rect 22500 4320 22564 4324
rect 22580 4380 22644 4384
rect 22580 4324 22584 4380
rect 22584 4324 22640 4380
rect 22640 4324 22644 4380
rect 22580 4320 22644 4324
rect 33034 4380 33098 4384
rect 33034 4324 33038 4380
rect 33038 4324 33094 4380
rect 33094 4324 33098 4380
rect 33034 4320 33098 4324
rect 33114 4380 33178 4384
rect 33114 4324 33118 4380
rect 33118 4324 33174 4380
rect 33174 4324 33178 4380
rect 33114 4320 33178 4324
rect 33194 4380 33258 4384
rect 33194 4324 33198 4380
rect 33198 4324 33254 4380
rect 33254 4324 33258 4380
rect 33194 4320 33258 4324
rect 33274 4380 33338 4384
rect 33274 4324 33278 4380
rect 33278 4324 33334 4380
rect 33334 4324 33338 4380
rect 33274 4320 33338 4324
rect 43728 4380 43792 4384
rect 43728 4324 43732 4380
rect 43732 4324 43788 4380
rect 43788 4324 43792 4380
rect 43728 4320 43792 4324
rect 43808 4380 43872 4384
rect 43808 4324 43812 4380
rect 43812 4324 43868 4380
rect 43868 4324 43872 4380
rect 43808 4320 43872 4324
rect 43888 4380 43952 4384
rect 43888 4324 43892 4380
rect 43892 4324 43948 4380
rect 43948 4324 43952 4380
rect 43888 4320 43952 4324
rect 43968 4380 44032 4384
rect 43968 4324 43972 4380
rect 43972 4324 44028 4380
rect 44028 4324 44032 4380
rect 43968 4320 44032 4324
rect 6299 3836 6363 3840
rect 6299 3780 6303 3836
rect 6303 3780 6359 3836
rect 6359 3780 6363 3836
rect 6299 3776 6363 3780
rect 6379 3836 6443 3840
rect 6379 3780 6383 3836
rect 6383 3780 6439 3836
rect 6439 3780 6443 3836
rect 6379 3776 6443 3780
rect 6459 3836 6523 3840
rect 6459 3780 6463 3836
rect 6463 3780 6519 3836
rect 6519 3780 6523 3836
rect 6459 3776 6523 3780
rect 6539 3836 6603 3840
rect 6539 3780 6543 3836
rect 6543 3780 6599 3836
rect 6599 3780 6603 3836
rect 6539 3776 6603 3780
rect 16993 3836 17057 3840
rect 16993 3780 16997 3836
rect 16997 3780 17053 3836
rect 17053 3780 17057 3836
rect 16993 3776 17057 3780
rect 17073 3836 17137 3840
rect 17073 3780 17077 3836
rect 17077 3780 17133 3836
rect 17133 3780 17137 3836
rect 17073 3776 17137 3780
rect 17153 3836 17217 3840
rect 17153 3780 17157 3836
rect 17157 3780 17213 3836
rect 17213 3780 17217 3836
rect 17153 3776 17217 3780
rect 17233 3836 17297 3840
rect 17233 3780 17237 3836
rect 17237 3780 17293 3836
rect 17293 3780 17297 3836
rect 17233 3776 17297 3780
rect 27687 3836 27751 3840
rect 27687 3780 27691 3836
rect 27691 3780 27747 3836
rect 27747 3780 27751 3836
rect 27687 3776 27751 3780
rect 27767 3836 27831 3840
rect 27767 3780 27771 3836
rect 27771 3780 27827 3836
rect 27827 3780 27831 3836
rect 27767 3776 27831 3780
rect 27847 3836 27911 3840
rect 27847 3780 27851 3836
rect 27851 3780 27907 3836
rect 27907 3780 27911 3836
rect 27847 3776 27911 3780
rect 27927 3836 27991 3840
rect 27927 3780 27931 3836
rect 27931 3780 27987 3836
rect 27987 3780 27991 3836
rect 27927 3776 27991 3780
rect 38381 3836 38445 3840
rect 38381 3780 38385 3836
rect 38385 3780 38441 3836
rect 38441 3780 38445 3836
rect 38381 3776 38445 3780
rect 38461 3836 38525 3840
rect 38461 3780 38465 3836
rect 38465 3780 38521 3836
rect 38521 3780 38525 3836
rect 38461 3776 38525 3780
rect 38541 3836 38605 3840
rect 38541 3780 38545 3836
rect 38545 3780 38601 3836
rect 38601 3780 38605 3836
rect 38541 3776 38605 3780
rect 38621 3836 38685 3840
rect 38621 3780 38625 3836
rect 38625 3780 38681 3836
rect 38681 3780 38685 3836
rect 38621 3776 38685 3780
rect 11646 3292 11710 3296
rect 11646 3236 11650 3292
rect 11650 3236 11706 3292
rect 11706 3236 11710 3292
rect 11646 3232 11710 3236
rect 11726 3292 11790 3296
rect 11726 3236 11730 3292
rect 11730 3236 11786 3292
rect 11786 3236 11790 3292
rect 11726 3232 11790 3236
rect 11806 3292 11870 3296
rect 11806 3236 11810 3292
rect 11810 3236 11866 3292
rect 11866 3236 11870 3292
rect 11806 3232 11870 3236
rect 11886 3292 11950 3296
rect 11886 3236 11890 3292
rect 11890 3236 11946 3292
rect 11946 3236 11950 3292
rect 11886 3232 11950 3236
rect 22340 3292 22404 3296
rect 22340 3236 22344 3292
rect 22344 3236 22400 3292
rect 22400 3236 22404 3292
rect 22340 3232 22404 3236
rect 22420 3292 22484 3296
rect 22420 3236 22424 3292
rect 22424 3236 22480 3292
rect 22480 3236 22484 3292
rect 22420 3232 22484 3236
rect 22500 3292 22564 3296
rect 22500 3236 22504 3292
rect 22504 3236 22560 3292
rect 22560 3236 22564 3292
rect 22500 3232 22564 3236
rect 22580 3292 22644 3296
rect 22580 3236 22584 3292
rect 22584 3236 22640 3292
rect 22640 3236 22644 3292
rect 22580 3232 22644 3236
rect 33034 3292 33098 3296
rect 33034 3236 33038 3292
rect 33038 3236 33094 3292
rect 33094 3236 33098 3292
rect 33034 3232 33098 3236
rect 33114 3292 33178 3296
rect 33114 3236 33118 3292
rect 33118 3236 33174 3292
rect 33174 3236 33178 3292
rect 33114 3232 33178 3236
rect 33194 3292 33258 3296
rect 33194 3236 33198 3292
rect 33198 3236 33254 3292
rect 33254 3236 33258 3292
rect 33194 3232 33258 3236
rect 33274 3292 33338 3296
rect 33274 3236 33278 3292
rect 33278 3236 33334 3292
rect 33334 3236 33338 3292
rect 33274 3232 33338 3236
rect 43728 3292 43792 3296
rect 43728 3236 43732 3292
rect 43732 3236 43788 3292
rect 43788 3236 43792 3292
rect 43728 3232 43792 3236
rect 43808 3292 43872 3296
rect 43808 3236 43812 3292
rect 43812 3236 43868 3292
rect 43868 3236 43872 3292
rect 43808 3232 43872 3236
rect 43888 3292 43952 3296
rect 43888 3236 43892 3292
rect 43892 3236 43948 3292
rect 43948 3236 43952 3292
rect 43888 3232 43952 3236
rect 43968 3292 44032 3296
rect 43968 3236 43972 3292
rect 43972 3236 44028 3292
rect 44028 3236 44032 3292
rect 43968 3232 44032 3236
rect 6299 2748 6363 2752
rect 6299 2692 6303 2748
rect 6303 2692 6359 2748
rect 6359 2692 6363 2748
rect 6299 2688 6363 2692
rect 6379 2748 6443 2752
rect 6379 2692 6383 2748
rect 6383 2692 6439 2748
rect 6439 2692 6443 2748
rect 6379 2688 6443 2692
rect 6459 2748 6523 2752
rect 6459 2692 6463 2748
rect 6463 2692 6519 2748
rect 6519 2692 6523 2748
rect 6459 2688 6523 2692
rect 6539 2748 6603 2752
rect 6539 2692 6543 2748
rect 6543 2692 6599 2748
rect 6599 2692 6603 2748
rect 6539 2688 6603 2692
rect 16993 2748 17057 2752
rect 16993 2692 16997 2748
rect 16997 2692 17053 2748
rect 17053 2692 17057 2748
rect 16993 2688 17057 2692
rect 17073 2748 17137 2752
rect 17073 2692 17077 2748
rect 17077 2692 17133 2748
rect 17133 2692 17137 2748
rect 17073 2688 17137 2692
rect 17153 2748 17217 2752
rect 17153 2692 17157 2748
rect 17157 2692 17213 2748
rect 17213 2692 17217 2748
rect 17153 2688 17217 2692
rect 17233 2748 17297 2752
rect 17233 2692 17237 2748
rect 17237 2692 17293 2748
rect 17293 2692 17297 2748
rect 17233 2688 17297 2692
rect 30236 2756 30300 2820
rect 36124 2756 36188 2820
rect 27687 2748 27751 2752
rect 27687 2692 27691 2748
rect 27691 2692 27747 2748
rect 27747 2692 27751 2748
rect 27687 2688 27751 2692
rect 27767 2748 27831 2752
rect 27767 2692 27771 2748
rect 27771 2692 27827 2748
rect 27827 2692 27831 2748
rect 27767 2688 27831 2692
rect 27847 2748 27911 2752
rect 27847 2692 27851 2748
rect 27851 2692 27907 2748
rect 27907 2692 27911 2748
rect 27847 2688 27911 2692
rect 27927 2748 27991 2752
rect 27927 2692 27931 2748
rect 27931 2692 27987 2748
rect 27987 2692 27991 2748
rect 27927 2688 27991 2692
rect 38381 2748 38445 2752
rect 38381 2692 38385 2748
rect 38385 2692 38441 2748
rect 38441 2692 38445 2748
rect 38381 2688 38445 2692
rect 38461 2748 38525 2752
rect 38461 2692 38465 2748
rect 38465 2692 38521 2748
rect 38521 2692 38525 2748
rect 38461 2688 38525 2692
rect 38541 2748 38605 2752
rect 38541 2692 38545 2748
rect 38545 2692 38601 2748
rect 38601 2692 38605 2748
rect 38541 2688 38605 2692
rect 38621 2748 38685 2752
rect 38621 2692 38625 2748
rect 38625 2692 38681 2748
rect 38681 2692 38685 2748
rect 38621 2688 38685 2692
rect 36860 2620 36924 2684
rect 11646 2204 11710 2208
rect 11646 2148 11650 2204
rect 11650 2148 11706 2204
rect 11706 2148 11710 2204
rect 11646 2144 11710 2148
rect 11726 2204 11790 2208
rect 11726 2148 11730 2204
rect 11730 2148 11786 2204
rect 11786 2148 11790 2204
rect 11726 2144 11790 2148
rect 11806 2204 11870 2208
rect 11806 2148 11810 2204
rect 11810 2148 11866 2204
rect 11866 2148 11870 2204
rect 11806 2144 11870 2148
rect 11886 2204 11950 2208
rect 11886 2148 11890 2204
rect 11890 2148 11946 2204
rect 11946 2148 11950 2204
rect 11886 2144 11950 2148
rect 22340 2204 22404 2208
rect 22340 2148 22344 2204
rect 22344 2148 22400 2204
rect 22400 2148 22404 2204
rect 22340 2144 22404 2148
rect 22420 2204 22484 2208
rect 22420 2148 22424 2204
rect 22424 2148 22480 2204
rect 22480 2148 22484 2204
rect 22420 2144 22484 2148
rect 22500 2204 22564 2208
rect 22500 2148 22504 2204
rect 22504 2148 22560 2204
rect 22560 2148 22564 2204
rect 22500 2144 22564 2148
rect 22580 2204 22644 2208
rect 22580 2148 22584 2204
rect 22584 2148 22640 2204
rect 22640 2148 22644 2204
rect 22580 2144 22644 2148
rect 33034 2204 33098 2208
rect 33034 2148 33038 2204
rect 33038 2148 33094 2204
rect 33094 2148 33098 2204
rect 33034 2144 33098 2148
rect 33114 2204 33178 2208
rect 33114 2148 33118 2204
rect 33118 2148 33174 2204
rect 33174 2148 33178 2204
rect 33114 2144 33178 2148
rect 33194 2204 33258 2208
rect 33194 2148 33198 2204
rect 33198 2148 33254 2204
rect 33254 2148 33258 2204
rect 33194 2144 33258 2148
rect 33274 2204 33338 2208
rect 33274 2148 33278 2204
rect 33278 2148 33334 2204
rect 33334 2148 33338 2204
rect 33274 2144 33338 2148
rect 43728 2204 43792 2208
rect 43728 2148 43732 2204
rect 43732 2148 43788 2204
rect 43788 2148 43792 2204
rect 43728 2144 43792 2148
rect 43808 2204 43872 2208
rect 43808 2148 43812 2204
rect 43812 2148 43868 2204
rect 43868 2148 43872 2204
rect 43808 2144 43872 2148
rect 43888 2204 43952 2208
rect 43888 2148 43892 2204
rect 43892 2148 43948 2204
rect 43948 2148 43952 2204
rect 43888 2144 43952 2148
rect 43968 2204 44032 2208
rect 43968 2148 43972 2204
rect 43972 2148 44028 2204
rect 44028 2148 44032 2204
rect 43968 2144 44032 2148
rect 30236 1260 30300 1324
rect 36124 852 36188 916
<< metal4 >>
rect 6291 7104 6611 7664
rect 6291 7040 6299 7104
rect 6363 7040 6379 7104
rect 6443 7040 6459 7104
rect 6523 7040 6539 7104
rect 6603 7040 6611 7104
rect 6291 6016 6611 7040
rect 6291 5952 6299 6016
rect 6363 5952 6379 6016
rect 6443 5952 6459 6016
rect 6523 5952 6539 6016
rect 6603 5952 6611 6016
rect 6291 4928 6611 5952
rect 6291 4864 6299 4928
rect 6363 4864 6379 4928
rect 6443 4864 6459 4928
rect 6523 4864 6539 4928
rect 6603 4864 6611 4928
rect 6291 3840 6611 4864
rect 6291 3776 6299 3840
rect 6363 3776 6379 3840
rect 6443 3776 6459 3840
rect 6523 3776 6539 3840
rect 6603 3776 6611 3840
rect 6291 2752 6611 3776
rect 6291 2688 6299 2752
rect 6363 2688 6379 2752
rect 6443 2688 6459 2752
rect 6523 2688 6539 2752
rect 6603 2688 6611 2752
rect 6291 2128 6611 2688
rect 11638 7648 11958 7664
rect 11638 7584 11646 7648
rect 11710 7584 11726 7648
rect 11790 7584 11806 7648
rect 11870 7584 11886 7648
rect 11950 7584 11958 7648
rect 11638 6560 11958 7584
rect 11638 6496 11646 6560
rect 11710 6496 11726 6560
rect 11790 6496 11806 6560
rect 11870 6496 11886 6560
rect 11950 6496 11958 6560
rect 11638 5472 11958 6496
rect 11638 5408 11646 5472
rect 11710 5408 11726 5472
rect 11790 5408 11806 5472
rect 11870 5408 11886 5472
rect 11950 5408 11958 5472
rect 11638 4384 11958 5408
rect 11638 4320 11646 4384
rect 11710 4320 11726 4384
rect 11790 4320 11806 4384
rect 11870 4320 11886 4384
rect 11950 4320 11958 4384
rect 11638 3296 11958 4320
rect 11638 3232 11646 3296
rect 11710 3232 11726 3296
rect 11790 3232 11806 3296
rect 11870 3232 11886 3296
rect 11950 3232 11958 3296
rect 11638 2208 11958 3232
rect 11638 2144 11646 2208
rect 11710 2144 11726 2208
rect 11790 2144 11806 2208
rect 11870 2144 11886 2208
rect 11950 2144 11958 2208
rect 11638 2128 11958 2144
rect 16985 7104 17305 7664
rect 16985 7040 16993 7104
rect 17057 7040 17073 7104
rect 17137 7040 17153 7104
rect 17217 7040 17233 7104
rect 17297 7040 17305 7104
rect 16985 6016 17305 7040
rect 16985 5952 16993 6016
rect 17057 5952 17073 6016
rect 17137 5952 17153 6016
rect 17217 5952 17233 6016
rect 17297 5952 17305 6016
rect 16985 4928 17305 5952
rect 16985 4864 16993 4928
rect 17057 4864 17073 4928
rect 17137 4864 17153 4928
rect 17217 4864 17233 4928
rect 17297 4864 17305 4928
rect 16985 3840 17305 4864
rect 16985 3776 16993 3840
rect 17057 3776 17073 3840
rect 17137 3776 17153 3840
rect 17217 3776 17233 3840
rect 17297 3776 17305 3840
rect 16985 2752 17305 3776
rect 16985 2688 16993 2752
rect 17057 2688 17073 2752
rect 17137 2688 17153 2752
rect 17217 2688 17233 2752
rect 17297 2688 17305 2752
rect 16985 2128 17305 2688
rect 22332 7648 22652 7664
rect 22332 7584 22340 7648
rect 22404 7584 22420 7648
rect 22484 7584 22500 7648
rect 22564 7584 22580 7648
rect 22644 7584 22652 7648
rect 22332 6560 22652 7584
rect 22332 6496 22340 6560
rect 22404 6496 22420 6560
rect 22484 6496 22500 6560
rect 22564 6496 22580 6560
rect 22644 6496 22652 6560
rect 22332 5472 22652 6496
rect 22332 5408 22340 5472
rect 22404 5408 22420 5472
rect 22484 5408 22500 5472
rect 22564 5408 22580 5472
rect 22644 5408 22652 5472
rect 22332 4384 22652 5408
rect 22332 4320 22340 4384
rect 22404 4320 22420 4384
rect 22484 4320 22500 4384
rect 22564 4320 22580 4384
rect 22644 4320 22652 4384
rect 22332 3296 22652 4320
rect 22332 3232 22340 3296
rect 22404 3232 22420 3296
rect 22484 3232 22500 3296
rect 22564 3232 22580 3296
rect 22644 3232 22652 3296
rect 22332 2208 22652 3232
rect 22332 2144 22340 2208
rect 22404 2144 22420 2208
rect 22484 2144 22500 2208
rect 22564 2144 22580 2208
rect 22644 2144 22652 2208
rect 22332 2128 22652 2144
rect 27679 7104 27999 7664
rect 27679 7040 27687 7104
rect 27751 7040 27767 7104
rect 27831 7040 27847 7104
rect 27911 7040 27927 7104
rect 27991 7040 27999 7104
rect 27679 6016 27999 7040
rect 27679 5952 27687 6016
rect 27751 5952 27767 6016
rect 27831 5952 27847 6016
rect 27911 5952 27927 6016
rect 27991 5952 27999 6016
rect 27679 4928 27999 5952
rect 27679 4864 27687 4928
rect 27751 4864 27767 4928
rect 27831 4864 27847 4928
rect 27911 4864 27927 4928
rect 27991 4864 27999 4928
rect 27679 3840 27999 4864
rect 27679 3776 27687 3840
rect 27751 3776 27767 3840
rect 27831 3776 27847 3840
rect 27911 3776 27927 3840
rect 27991 3776 27999 3840
rect 27679 2752 27999 3776
rect 33026 7648 33346 7664
rect 33026 7584 33034 7648
rect 33098 7584 33114 7648
rect 33178 7584 33194 7648
rect 33258 7584 33274 7648
rect 33338 7584 33346 7648
rect 33026 6560 33346 7584
rect 33026 6496 33034 6560
rect 33098 6496 33114 6560
rect 33178 6496 33194 6560
rect 33258 6496 33274 6560
rect 33338 6496 33346 6560
rect 33026 5472 33346 6496
rect 38373 7104 38693 7664
rect 38373 7040 38381 7104
rect 38445 7040 38461 7104
rect 38525 7040 38541 7104
rect 38605 7040 38621 7104
rect 38685 7040 38693 7104
rect 38373 6016 38693 7040
rect 38373 5952 38381 6016
rect 38445 5952 38461 6016
rect 38525 5952 38541 6016
rect 38605 5952 38621 6016
rect 38685 5952 38693 6016
rect 36859 5676 36925 5677
rect 36859 5612 36860 5676
rect 36924 5612 36925 5676
rect 36859 5611 36925 5612
rect 33026 5408 33034 5472
rect 33098 5408 33114 5472
rect 33178 5408 33194 5472
rect 33258 5408 33274 5472
rect 33338 5408 33346 5472
rect 33026 4384 33346 5408
rect 33026 4320 33034 4384
rect 33098 4320 33114 4384
rect 33178 4320 33194 4384
rect 33258 4320 33274 4384
rect 33338 4320 33346 4384
rect 33026 3296 33346 4320
rect 33026 3232 33034 3296
rect 33098 3232 33114 3296
rect 33178 3232 33194 3296
rect 33258 3232 33274 3296
rect 33338 3232 33346 3296
rect 30235 2820 30301 2821
rect 30235 2756 30236 2820
rect 30300 2756 30301 2820
rect 30235 2755 30301 2756
rect 27679 2688 27687 2752
rect 27751 2688 27767 2752
rect 27831 2688 27847 2752
rect 27911 2688 27927 2752
rect 27991 2688 27999 2752
rect 27679 2128 27999 2688
rect 30238 1325 30298 2755
rect 33026 2208 33346 3232
rect 36123 2820 36189 2821
rect 36123 2756 36124 2820
rect 36188 2756 36189 2820
rect 36123 2755 36189 2756
rect 33026 2144 33034 2208
rect 33098 2144 33114 2208
rect 33178 2144 33194 2208
rect 33258 2144 33274 2208
rect 33338 2144 33346 2208
rect 33026 2128 33346 2144
rect 30235 1324 30301 1325
rect 30235 1260 30236 1324
rect 30300 1260 30301 1324
rect 30235 1259 30301 1260
rect 36126 917 36186 2755
rect 36862 2685 36922 5611
rect 38373 4928 38693 5952
rect 38373 4864 38381 4928
rect 38445 4864 38461 4928
rect 38525 4864 38541 4928
rect 38605 4864 38621 4928
rect 38685 4864 38693 4928
rect 38373 3840 38693 4864
rect 38373 3776 38381 3840
rect 38445 3776 38461 3840
rect 38525 3776 38541 3840
rect 38605 3776 38621 3840
rect 38685 3776 38693 3840
rect 38373 2752 38693 3776
rect 38373 2688 38381 2752
rect 38445 2688 38461 2752
rect 38525 2688 38541 2752
rect 38605 2688 38621 2752
rect 38685 2688 38693 2752
rect 36859 2684 36925 2685
rect 36859 2620 36860 2684
rect 36924 2620 36925 2684
rect 36859 2619 36925 2620
rect 38373 2128 38693 2688
rect 43720 7648 44040 7664
rect 43720 7584 43728 7648
rect 43792 7584 43808 7648
rect 43872 7584 43888 7648
rect 43952 7584 43968 7648
rect 44032 7584 44040 7648
rect 43720 6560 44040 7584
rect 43720 6496 43728 6560
rect 43792 6496 43808 6560
rect 43872 6496 43888 6560
rect 43952 6496 43968 6560
rect 44032 6496 44040 6560
rect 43720 5472 44040 6496
rect 43720 5408 43728 5472
rect 43792 5408 43808 5472
rect 43872 5408 43888 5472
rect 43952 5408 43968 5472
rect 44032 5408 44040 5472
rect 43720 4384 44040 5408
rect 43720 4320 43728 4384
rect 43792 4320 43808 4384
rect 43872 4320 43888 4384
rect 43952 4320 43968 4384
rect 44032 4320 44040 4384
rect 43720 3296 44040 4320
rect 43720 3232 43728 3296
rect 43792 3232 43808 3296
rect 43872 3232 43888 3296
rect 43952 3232 43968 3296
rect 44032 3232 44040 3296
rect 43720 2208 44040 3232
rect 43720 2144 43728 2208
rect 43792 2144 43808 2208
rect 43872 2144 43888 2208
rect 43952 2144 43968 2208
rect 44032 2144 44040 2208
rect 43720 2128 44040 2144
rect 36123 916 36189 917
rect 36123 852 36124 916
rect 36188 852 36189 916
rect 36123 851 36189 852
use sky130_fd_sc_hd__clkbuf_1  _00_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _01_
timestamp 1688980957
transform 1 0 20976 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp 1688980957
transform 1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1688980957
transform 1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1688980957
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1688980957
transform 1 0 37904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1688980957
transform 1 0 38088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 40388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 41216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 42780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1688980957
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1688980957
transform 1 0 23736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1688980957
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1688980957
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1688980957
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1688980957
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1688980957
transform 1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1688980957
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1688980957
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1688980957
transform 1 0 25760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1688980957
transform 1 0 26036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1688980957
transform 1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1688980957
transform 1 0 26864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1688980957
transform 1 0 27232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1688980957
transform 1 0 27784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1688980957
transform 1 0 28060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1688980957
transform 1 0 28336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1688980957
transform 1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _49_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _50_
timestamp 1688980957
transform 1 0 18952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _51_
timestamp 1688980957
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _52_
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _53_
timestamp 1688980957
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _54_
timestamp 1688980957
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _55_
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _56_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _57_
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _58_
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _59_
timestamp 1688980957
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _60_
timestamp 1688980957
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _61_
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _62_
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _63_
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _64_
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _65_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _66_
timestamp 1688980957
transform -1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _67_
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _68_
timestamp 1688980957
transform 1 0 34868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _69_
timestamp 1688980957
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _70_
timestamp 1688980957
transform 1 0 35236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1688980957
transform -1 0 16652 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform -1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 32292 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_144 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_148
timestamp 1688980957
transform 1 0 14720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1688980957
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_439
timestamp 1688980957
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_447
timestamp 1688980957
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_449 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_456 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43056 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_90
timestamp 1688980957
transform 1 0 9384 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_102
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_140
timestamp 1688980957
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_341
timestamp 1688980957
transform 1 0 32476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_384
timestamp 1688980957
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_174 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_180
timestamp 1688980957
transform 1 0 17664 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_188
timestamp 1688980957
transform 1 0 18400 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp 1688980957
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_208
timestamp 1688980957
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_230
timestamp 1688980957
transform 1 0 22264 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_235
timestamp 1688980957
transform 1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_244
timestamp 1688980957
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_259
timestamp 1688980957
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_283
timestamp 1688980957
transform 1 0 27140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_287
timestamp 1688980957
transform 1 0 27508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_302
timestamp 1688980957
transform 1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_355
timestamp 1688980957
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_461
timestamp 1688980957
transform 1 0 43516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_461
timestamp 1688980957
transform 1 0 43516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_161
timestamp 1688980957
transform 1 0 15916 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_164
timestamp 1688980957
transform 1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_169
timestamp 1688980957
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_181
timestamp 1688980957
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_193
timestamp 1688980957
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_257
timestamp 1688980957
transform 1 0 24748 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_261
timestamp 1688980957
transform 1 0 25116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_273
timestamp 1688980957
transform 1 0 26220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_285
timestamp 1688980957
transform 1 0 27324 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_297
timestamp 1688980957
transform 1 0 28428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_305
timestamp 1688980957
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_461
timestamp 1688980957
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_239
timestamp 1688980957
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_461
timestamp 1688980957
transform 1 0 43516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_21
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_35
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_47
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_78
timestamp 1688980957
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_85
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_101
timestamp 1688980957
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 1688980957
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_117
timestamp 1688980957
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_124
timestamp 1688980957
transform 1 0 12512 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_136
timestamp 1688980957
transform 1 0 13616 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_147
timestamp 1688980957
transform 1 0 14628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_159
timestamp 1688980957
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_175
timestamp 1688980957
transform 1 0 17204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_197
timestamp 1688980957
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_209
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_219
timestamp 1688980957
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_233
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_248
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_253
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_262
timestamp 1688980957
transform 1 0 25208 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_274
timestamp 1688980957
transform 1 0 26312 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_290
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_309
timestamp 1688980957
transform 1 0 29532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_321
timestamp 1688980957
transform 1 0 30636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_331
timestamp 1688980957
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_345
timestamp 1688980957
transform 1 0 32844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_354
timestamp 1688980957
transform 1 0 33672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_362
timestamp 1688980957
transform 1 0 34408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_365
timestamp 1688980957
transform 1 0 34684 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_377
timestamp 1688980957
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_389
timestamp 1688980957
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_403
timestamp 1688980957
transform 1 0 38180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_415
timestamp 1688980957
transform 1 0 39284 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_419
timestamp 1688980957
transform 1 0 39652 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_427
timestamp 1688980957
transform 1 0 40388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_439
timestamp 1688980957
transform 1 0 41492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_446
timestamp 1688980957
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_455
timestamp 1688980957
transform 1 0 42964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 36524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 38640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 38916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 37812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 38916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 39192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 36800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 35880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 38088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 17572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 18400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 19320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform 1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform 1 0 16744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform 1 0 17296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 24656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 28888 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 31004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 33120 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 35236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 37352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 39836 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 41584 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 43056 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 11960 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 18308 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 20424 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 23368 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 23184 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 24932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 24564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 20608 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 22080 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 22080 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 28612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 30084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 29716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 26036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 25668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 27508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 33764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 31188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 30820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 32660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 33764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 32660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal2 s 34150 0 34206 160 0 FreeSans 224 90 0 0 Ci
port 0 nsew signal input
flabel metal2 s 34426 0 34482 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 1 nsew signal input
flabel metal2 s 37186 0 37242 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 2 nsew signal input
flabel metal2 s 37462 0 37518 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 3 nsew signal input
flabel metal2 s 37738 0 37794 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 4 nsew signal input
flabel metal2 s 38014 0 38070 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 5 nsew signal input
flabel metal2 s 38290 0 38346 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 6 nsew signal input
flabel metal2 s 38566 0 38622 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 7 nsew signal input
flabel metal2 s 38842 0 38898 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 8 nsew signal input
flabel metal2 s 39118 0 39174 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 9 nsew signal input
flabel metal2 s 39394 0 39450 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 10 nsew signal input
flabel metal2 s 39670 0 39726 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 11 nsew signal input
flabel metal2 s 34702 0 34758 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 12 nsew signal input
flabel metal2 s 34978 0 35034 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 13 nsew signal input
flabel metal2 s 35254 0 35310 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 14 nsew signal input
flabel metal2 s 35530 0 35586 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 15 nsew signal input
flabel metal2 s 35806 0 35862 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 16 nsew signal input
flabel metal2 s 36082 0 36138 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 17 nsew signal input
flabel metal2 s 36358 0 36414 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 18 nsew signal input
flabel metal2 s 36634 0 36690 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 19 nsew signal input
flabel metal2 s 36910 0 36966 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 20 nsew signal input
flabel metal2 s 3422 9840 3478 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 21 nsew signal tristate
flabel metal2 s 24582 9840 24638 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 22 nsew signal tristate
flabel metal2 s 26698 9840 26754 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 23 nsew signal tristate
flabel metal2 s 28814 9840 28870 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 24 nsew signal tristate
flabel metal2 s 30930 9840 30986 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 25 nsew signal tristate
flabel metal2 s 33046 9840 33102 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 26 nsew signal tristate
flabel metal2 s 35162 9840 35218 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 27 nsew signal tristate
flabel metal2 s 37278 9840 37334 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 28 nsew signal tristate
flabel metal2 s 39394 9840 39450 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 29 nsew signal tristate
flabel metal2 s 41510 9840 41566 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 30 nsew signal tristate
flabel metal2 s 43626 9840 43682 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 31 nsew signal tristate
flabel metal2 s 5538 9840 5594 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 32 nsew signal tristate
flabel metal2 s 7654 9840 7710 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 33 nsew signal tristate
flabel metal2 s 9770 9840 9826 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 34 nsew signal tristate
flabel metal2 s 11886 9840 11942 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 35 nsew signal tristate
flabel metal2 s 14002 9840 14058 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 36 nsew signal tristate
flabel metal2 s 16118 9840 16174 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 37 nsew signal tristate
flabel metal2 s 18234 9840 18290 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 38 nsew signal tristate
flabel metal2 s 20350 9840 20406 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 39 nsew signal tristate
flabel metal2 s 22466 9840 22522 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 40 nsew signal tristate
flabel metal2 s 5170 0 5226 160 0 FreeSans 224 90 0 0 N1END[0]
port 41 nsew signal input
flabel metal2 s 5446 0 5502 160 0 FreeSans 224 90 0 0 N1END[1]
port 42 nsew signal input
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 N1END[2]
port 43 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 N1END[3]
port 44 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N2END[0]
port 45 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N2END[1]
port 46 nsew signal input
flabel metal2 s 9034 0 9090 160 0 FreeSans 224 90 0 0 N2END[2]
port 47 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 N2END[3]
port 48 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N2END[4]
port 49 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N2END[5]
port 50 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 N2END[6]
port 51 nsew signal input
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 N2END[7]
port 52 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N2MID[0]
port 53 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N2MID[1]
port 54 nsew signal input
flabel metal2 s 6826 0 6882 160 0 FreeSans 224 90 0 0 N2MID[2]
port 55 nsew signal input
flabel metal2 s 7102 0 7158 160 0 FreeSans 224 90 0 0 N2MID[3]
port 56 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N2MID[4]
port 57 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N2MID[5]
port 58 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 N2MID[6]
port 59 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 N2MID[7]
port 60 nsew signal input
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 N4END[0]
port 61 nsew signal input
flabel metal2 s 13450 0 13506 160 0 FreeSans 224 90 0 0 N4END[10]
port 62 nsew signal input
flabel metal2 s 13726 0 13782 160 0 FreeSans 224 90 0 0 N4END[11]
port 63 nsew signal input
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 N4END[12]
port 64 nsew signal input
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 N4END[13]
port 65 nsew signal input
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 N4END[14]
port 66 nsew signal input
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 N4END[15]
port 67 nsew signal input
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 N4END[1]
port 68 nsew signal input
flabel metal2 s 11242 0 11298 160 0 FreeSans 224 90 0 0 N4END[2]
port 69 nsew signal input
flabel metal2 s 11518 0 11574 160 0 FreeSans 224 90 0 0 N4END[3]
port 70 nsew signal input
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 N4END[4]
port 71 nsew signal input
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 N4END[5]
port 72 nsew signal input
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 N4END[6]
port 73 nsew signal input
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 N4END[7]
port 74 nsew signal input
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 N4END[8]
port 75 nsew signal input
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 N4END[9]
port 76 nsew signal input
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 NN4END[0]
port 77 nsew signal input
flabel metal2 s 17866 0 17922 160 0 FreeSans 224 90 0 0 NN4END[10]
port 78 nsew signal input
flabel metal2 s 18142 0 18198 160 0 FreeSans 224 90 0 0 NN4END[11]
port 79 nsew signal input
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 NN4END[12]
port 80 nsew signal input
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 NN4END[13]
port 81 nsew signal input
flabel metal2 s 18970 0 19026 160 0 FreeSans 224 90 0 0 NN4END[14]
port 82 nsew signal input
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 NN4END[15]
port 83 nsew signal input
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 NN4END[1]
port 84 nsew signal input
flabel metal2 s 15658 0 15714 160 0 FreeSans 224 90 0 0 NN4END[2]
port 85 nsew signal input
flabel metal2 s 15934 0 15990 160 0 FreeSans 224 90 0 0 NN4END[3]
port 86 nsew signal input
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 NN4END[4]
port 87 nsew signal input
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 NN4END[5]
port 88 nsew signal input
flabel metal2 s 16762 0 16818 160 0 FreeSans 224 90 0 0 NN4END[6]
port 89 nsew signal input
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 NN4END[7]
port 90 nsew signal input
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 NN4END[8]
port 91 nsew signal input
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 NN4END[9]
port 92 nsew signal input
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 93 nsew signal tristate
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 94 nsew signal tristate
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 95 nsew signal tristate
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 96 nsew signal tristate
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 97 nsew signal tristate
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 98 nsew signal tristate
flabel metal2 s 23386 0 23442 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 99 nsew signal tristate
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 100 nsew signal tristate
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 101 nsew signal tristate
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 102 nsew signal tristate
flabel metal2 s 24490 0 24546 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 103 nsew signal tristate
flabel metal2 s 24766 0 24822 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 104 nsew signal tristate
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 105 nsew signal tristate
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 106 nsew signal tristate
flabel metal2 s 21178 0 21234 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 107 nsew signal tristate
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 108 nsew signal tristate
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 109 nsew signal tristate
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 110 nsew signal tristate
flabel metal2 s 22282 0 22338 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 111 nsew signal tristate
flabel metal2 s 22558 0 22614 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 112 nsew signal tristate
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 113 nsew signal tristate
flabel metal2 s 27802 0 27858 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 114 nsew signal tristate
flabel metal2 s 28078 0 28134 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 115 nsew signal tristate
flabel metal2 s 28354 0 28410 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 116 nsew signal tristate
flabel metal2 s 28630 0 28686 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 117 nsew signal tristate
flabel metal2 s 28906 0 28962 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 118 nsew signal tristate
flabel metal2 s 29182 0 29238 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 119 nsew signal tristate
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 120 nsew signal tristate
flabel metal2 s 25594 0 25650 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 121 nsew signal tristate
flabel metal2 s 25870 0 25926 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 122 nsew signal tristate
flabel metal2 s 26146 0 26202 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 123 nsew signal tristate
flabel metal2 s 26422 0 26478 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 124 nsew signal tristate
flabel metal2 s 26698 0 26754 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 125 nsew signal tristate
flabel metal2 s 26974 0 27030 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 126 nsew signal tristate
flabel metal2 s 27250 0 27306 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 127 nsew signal tristate
flabel metal2 s 27526 0 27582 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 128 nsew signal tristate
flabel metal2 s 29458 0 29514 160 0 FreeSans 224 90 0 0 SS4BEG[0]
port 129 nsew signal tristate
flabel metal2 s 32218 0 32274 160 0 FreeSans 224 90 0 0 SS4BEG[10]
port 130 nsew signal tristate
flabel metal2 s 32494 0 32550 160 0 FreeSans 224 90 0 0 SS4BEG[11]
port 131 nsew signal tristate
flabel metal2 s 32770 0 32826 160 0 FreeSans 224 90 0 0 SS4BEG[12]
port 132 nsew signal tristate
flabel metal2 s 33046 0 33102 160 0 FreeSans 224 90 0 0 SS4BEG[13]
port 133 nsew signal tristate
flabel metal2 s 33322 0 33378 160 0 FreeSans 224 90 0 0 SS4BEG[14]
port 134 nsew signal tristate
flabel metal2 s 33598 0 33654 160 0 FreeSans 224 90 0 0 SS4BEG[15]
port 135 nsew signal tristate
flabel metal2 s 29734 0 29790 160 0 FreeSans 224 90 0 0 SS4BEG[1]
port 136 nsew signal tristate
flabel metal2 s 30010 0 30066 160 0 FreeSans 224 90 0 0 SS4BEG[2]
port 137 nsew signal tristate
flabel metal2 s 30286 0 30342 160 0 FreeSans 224 90 0 0 SS4BEG[3]
port 138 nsew signal tristate
flabel metal2 s 30562 0 30618 160 0 FreeSans 224 90 0 0 SS4BEG[4]
port 139 nsew signal tristate
flabel metal2 s 30838 0 30894 160 0 FreeSans 224 90 0 0 SS4BEG[5]
port 140 nsew signal tristate
flabel metal2 s 31114 0 31170 160 0 FreeSans 224 90 0 0 SS4BEG[6]
port 141 nsew signal tristate
flabel metal2 s 31390 0 31446 160 0 FreeSans 224 90 0 0 SS4BEG[7]
port 142 nsew signal tristate
flabel metal2 s 31666 0 31722 160 0 FreeSans 224 90 0 0 SS4BEG[8]
port 143 nsew signal tristate
flabel metal2 s 31942 0 31998 160 0 FreeSans 224 90 0 0 SS4BEG[9]
port 144 nsew signal tristate
flabel metal2 s 33874 0 33930 160 0 FreeSans 224 90 0 0 UserCLK
port 145 nsew signal input
flabel metal2 s 1306 9840 1362 10000 0 FreeSans 224 90 0 0 UserCLKo
port 146 nsew signal tristate
flabel metal4 s 6291 2128 6611 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 16985 2128 17305 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 27679 2128 27999 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 38373 2128 38693 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 11638 2128 11958 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 22332 2128 22652 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 33026 2128 33346 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 43720 2128 44040 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
rlabel metal1 22494 7072 22494 7072 0 vccd1
rlabel via1 22572 7616 22572 7616 0 vssd1
rlabel metal2 36570 1972 36570 1972 0 FrameStrobe[0]
rlabel metal2 37214 1452 37214 1452 0 FrameStrobe[10]
rlabel metal2 37490 687 37490 687 0 FrameStrobe[11]
rlabel metal2 37766 1554 37766 1554 0 FrameStrobe[12]
rlabel metal2 38042 738 38042 738 0 FrameStrobe[13]
rlabel metal2 38318 687 38318 687 0 FrameStrobe[14]
rlabel metal2 38594 772 38594 772 0 FrameStrobe[15]
rlabel metal2 38870 1554 38870 1554 0 FrameStrobe[16]
rlabel metal2 39146 823 39146 823 0 FrameStrobe[17]
rlabel metal2 39422 738 39422 738 0 FrameStrobe[18]
rlabel metal2 39698 143 39698 143 0 FrameStrobe[19]
rlabel metal2 34730 1520 34730 1520 0 FrameStrobe[1]
rlabel metal2 37030 2074 37030 2074 0 FrameStrobe[2]
rlabel metal1 36110 3060 36110 3060 0 FrameStrobe[3]
rlabel metal1 37490 1496 37490 1496 0 FrameStrobe[4]
rlabel metal1 36202 2992 36202 2992 0 FrameStrobe[5]
rlabel metal2 36110 687 36110 687 0 FrameStrobe[6]
rlabel metal2 36485 68 36485 68 0 FrameStrobe[7]
rlabel metal2 36761 68 36761 68 0 FrameStrobe[8]
rlabel metal2 37037 68 37037 68 0 FrameStrobe[9]
rlabel metal2 3450 9785 3450 9785 0 FrameStrobe_O[0]
rlabel metal2 24610 8629 24610 8629 0 FrameStrobe_O[10]
rlabel metal2 26726 8680 26726 8680 0 FrameStrobe_O[11]
rlabel metal2 28842 8629 28842 8629 0 FrameStrobe_O[12]
rlabel metal2 30958 8680 30958 8680 0 FrameStrobe_O[13]
rlabel metal2 33074 9173 33074 9173 0 FrameStrobe_O[14]
rlabel metal2 35190 8680 35190 8680 0 FrameStrobe_O[15]
rlabel metal2 37306 8680 37306 8680 0 FrameStrobe_O[16]
rlabel metal2 39422 9785 39422 9785 0 FrameStrobe_O[17]
rlabel metal2 41538 8680 41538 8680 0 FrameStrobe_O[18]
rlabel metal1 43562 7514 43562 7514 0 FrameStrobe_O[19]
rlabel metal2 5566 8680 5566 8680 0 FrameStrobe_O[1]
rlabel metal2 7682 8680 7682 8680 0 FrameStrobe_O[2]
rlabel metal2 9798 8680 9798 8680 0 FrameStrobe_O[3]
rlabel metal2 11914 9785 11914 9785 0 FrameStrobe_O[4]
rlabel metal2 14030 8680 14030 8680 0 FrameStrobe_O[5]
rlabel metal2 16146 9785 16146 9785 0 FrameStrobe_O[6]
rlabel metal2 18262 8510 18262 8510 0 FrameStrobe_O[7]
rlabel metal2 20378 9785 20378 9785 0 FrameStrobe_O[8]
rlabel metal2 22494 9785 22494 9785 0 FrameStrobe_O[9]
rlabel metal2 5198 1214 5198 1214 0 N1END[0]
rlabel metal2 5474 1214 5474 1214 0 N1END[1]
rlabel metal2 5750 1231 5750 1231 0 N1END[2]
rlabel metal2 6026 687 6026 687 0 N1END[3]
rlabel metal2 8510 1214 8510 1214 0 N2END[0]
rlabel metal2 8733 68 8733 68 0 N2END[1]
rlabel metal2 9115 68 9115 68 0 N2END[2]
rlabel metal2 9338 806 9338 806 0 N2END[3]
rlabel metal2 9614 1214 9614 1214 0 N2END[4]
rlabel metal2 9890 1282 9890 1282 0 N2END[5]
rlabel metal2 10166 1214 10166 1214 0 N2END[6]
rlabel metal2 10442 1282 10442 1282 0 N2END[7]
rlabel metal2 6302 738 6302 738 0 N2MID[0]
rlabel metal2 6479 68 6479 68 0 N2MID[1]
rlabel metal2 6854 687 6854 687 0 N2MID[2]
rlabel metal1 6670 2380 6670 2380 0 N2MID[3]
rlabel metal2 7353 68 7353 68 0 N2MID[4]
rlabel metal2 7583 68 7583 68 0 N2MID[5]
rlabel metal2 7859 68 7859 68 0 N2MID[6]
rlabel metal2 8135 68 8135 68 0 N2MID[7]
rlabel metal2 10718 1214 10718 1214 0 N4END[0]
rlabel metal2 13478 1214 13478 1214 0 N4END[10]
rlabel metal2 13754 1248 13754 1248 0 N4END[11]
rlabel metal1 13892 3026 13892 3026 0 N4END[12]
rlabel metal2 14306 1421 14306 1421 0 N4END[13]
rlabel metal2 14635 68 14635 68 0 N4END[14]
rlabel metal2 14911 68 14911 68 0 N4END[15]
rlabel metal2 10994 1282 10994 1282 0 N4END[1]
rlabel metal2 11270 1214 11270 1214 0 N4END[2]
rlabel metal2 11546 1299 11546 1299 0 N4END[3]
rlabel metal2 11822 738 11822 738 0 N4END[4]
rlabel metal2 12098 1214 12098 1214 0 N4END[5]
rlabel metal2 12374 1180 12374 1180 0 N4END[6]
rlabel metal2 12650 1214 12650 1214 0 N4END[7]
rlabel metal2 12926 1282 12926 1282 0 N4END[8]
rlabel metal2 13202 738 13202 738 0 N4END[9]
rlabel metal2 15081 68 15081 68 0 NN4END[0]
rlabel metal2 17848 2822 17848 2822 0 NN4END[10]
rlabel metal2 18170 636 18170 636 0 NN4END[11]
rlabel metal1 18584 3502 18584 3502 0 NN4END[12]
rlabel metal2 18722 959 18722 959 0 NN4END[13]
rlabel metal2 18998 1027 18998 1027 0 NN4END[14]
rlabel metal1 19412 3502 19412 3502 0 NN4END[15]
rlabel metal2 15410 1554 15410 1554 0 NN4END[1]
rlabel metal2 15686 1554 15686 1554 0 NN4END[2]
rlabel metal2 15962 1554 15962 1554 0 NN4END[3]
rlabel metal2 16238 1554 16238 1554 0 NN4END[4]
rlabel metal2 16514 1554 16514 1554 0 NN4END[5]
rlabel metal1 16928 3502 16928 3502 0 NN4END[6]
rlabel metal2 17066 823 17066 823 0 NN4END[7]
rlabel metal2 17395 68 17395 68 0 NN4END[8]
rlabel metal2 17572 2924 17572 2924 0 NN4END[9]
rlabel metal2 19550 1214 19550 1214 0 S1BEG[0]
rlabel metal2 19826 1486 19826 1486 0 S1BEG[1]
rlabel metal2 20201 68 20201 68 0 S1BEG[2]
rlabel metal2 20378 1214 20378 1214 0 S1BEG[3]
rlabel metal2 22862 1180 22862 1180 0 S2BEG[0]
rlabel metal1 23276 2822 23276 2822 0 S2BEG[1]
rlabel metal2 23414 755 23414 755 0 S2BEG[2]
rlabel metal2 23690 1180 23690 1180 0 S2BEG[3]
rlabel metal2 23966 619 23966 619 0 S2BEG[4]
rlabel metal2 24341 68 24341 68 0 S2BEG[5]
rlabel metal1 24656 2822 24656 2822 0 S2BEG[6]
rlabel metal2 24794 1350 24794 1350 0 S2BEG[7]
rlabel metal1 20746 2822 20746 2822 0 S2BEGb[0]
rlabel metal2 20831 68 20831 68 0 S2BEGb[1]
rlabel metal2 21305 68 21305 68 0 S2BEGb[2]
rlabel metal2 21482 1214 21482 1214 0 S2BEGb[3]
rlabel metal2 21705 68 21705 68 0 S2BEGb[4]
rlabel metal2 22034 1486 22034 1486 0 S2BEGb[5]
rlabel metal2 22257 68 22257 68 0 S2BEGb[6]
rlabel metal2 22685 68 22685 68 0 S2BEGb[7]
rlabel metal1 25208 2822 25208 2822 0 S4BEG[0]
rlabel metal2 27929 68 27929 68 0 S4BEG[10]
rlabel metal2 28205 68 28205 68 0 S4BEG[11]
rlabel metal2 28382 1180 28382 1180 0 S4BEG[12]
rlabel metal2 28757 68 28757 68 0 S4BEG[13]
rlabel metal2 28934 1316 28934 1316 0 S4BEG[14]
rlabel metal2 29348 2788 29348 2788 0 S4BEG[15]
rlabel metal2 25445 68 25445 68 0 S4BEG[1]
rlabel metal1 25760 2822 25760 2822 0 S4BEG[2]
rlabel metal2 25997 68 25997 68 0 S4BEG[3]
rlabel metal2 26174 755 26174 755 0 S4BEG[4]
rlabel metal2 26549 68 26549 68 0 S4BEG[5]
rlabel metal2 26825 68 26825 68 0 S4BEG[6]
rlabel metal1 27140 2890 27140 2890 0 S4BEG[7]
rlabel metal2 27377 68 27377 68 0 S4BEG[8]
rlabel metal1 27922 2890 27922 2890 0 S4BEG[9]
rlabel metal2 29585 68 29585 68 0 SS4BEG[0]
rlabel metal2 32345 68 32345 68 0 SS4BEG[10]
rlabel metal2 32522 1486 32522 1486 0 SS4BEG[11]
rlabel metal2 32798 1724 32798 1724 0 SS4BEG[12]
rlabel metal2 33021 68 33021 68 0 SS4BEG[13]
rlabel metal2 33403 68 33403 68 0 SS4BEG[14]
rlabel metal2 33626 1486 33626 1486 0 SS4BEG[15]
rlabel metal1 29900 2890 29900 2890 0 SS4BEG[1]
rlabel metal2 30137 68 30137 68 0 SS4BEG[2]
rlabel metal1 30682 2890 30682 2890 0 SS4BEG[3]
rlabel metal1 31096 3162 31096 3162 0 SS4BEG[4]
rlabel metal1 32890 2584 32890 2584 0 SS4BEG[5]
rlabel metal1 32683 2482 32683 2482 0 SS4BEG[6]
rlabel metal2 31517 68 31517 68 0 SS4BEG[7]
rlabel via1 31878 1445 31878 1445 0 SS4BEG[8]
rlabel metal2 31970 1486 31970 1486 0 SS4BEG[9]
rlabel metal2 34001 68 34001 68 0 UserCLK
rlabel metal2 1334 8680 1334 8680 0 UserCLKo
rlabel metal2 36754 4794 36754 4794 0 net1
rlabel metal1 41446 2448 41446 2448 0 net10
rlabel metal1 23322 2482 23322 2482 0 net100
rlabel metal1 23690 2414 23690 2414 0 net101
rlabel metal1 24242 2414 24242 2414 0 net102
rlabel metal1 24978 2414 24978 2414 0 net103
rlabel metal1 24702 3128 24702 3128 0 net104
rlabel metal1 25300 2346 25300 2346 0 net105
rlabel metal1 20746 3128 20746 3128 0 net106
rlabel metal1 20194 2448 20194 2448 0 net107
rlabel metal1 21068 3094 21068 3094 0 net108
rlabel metal1 20838 2414 20838 2414 0 net109
rlabel metal1 43010 2482 43010 2482 0 net11
rlabel metal1 21252 2414 21252 2414 0 net110
rlabel metal1 21482 3128 21482 3128 0 net111
rlabel metal1 21758 3400 21758 3400 0 net112
rlabel metal2 22034 3264 22034 3264 0 net113
rlabel metal1 24932 3026 24932 3026 0 net114
rlabel metal1 28014 3434 28014 3434 0 net115
rlabel metal1 29118 2618 29118 2618 0 net116
rlabel metal1 29624 2414 29624 2414 0 net117
rlabel metal1 28704 3094 28704 3094 0 net118
rlabel metal1 30038 2414 30038 2414 0 net119
rlabel metal2 36018 2652 36018 2652 0 net12
rlabel metal1 29854 3128 29854 3128 0 net120
rlabel metal1 25944 2414 25944 2414 0 net121
rlabel metal1 26450 2618 26450 2618 0 net122
rlabel metal1 26358 3060 26358 3060 0 net123
rlabel metal1 26312 3706 26312 3706 0 net124
rlabel metal1 26910 3026 26910 3026 0 net125
rlabel metal1 26956 2346 26956 2346 0 net126
rlabel metal1 27646 3128 27646 3128 0 net127
rlabel metal1 28152 2414 28152 2414 0 net128
rlabel metal1 27876 3026 27876 3026 0 net129
rlabel metal1 36892 2618 36892 2618 0 net13
rlabel metal1 19458 2924 19458 2924 0 net130
rlabel metal2 16606 1683 16606 1683 0 net131
rlabel metal2 16146 1734 16146 1734 0 net132
rlabel metal2 15870 1700 15870 1700 0 net133
rlabel metal2 15594 1768 15594 1768 0 net134
rlabel metal2 15134 1802 15134 1802 0 net135
rlabel metal1 33948 3094 33948 3094 0 net136
rlabel metal2 19182 3451 19182 3451 0 net137
rlabel metal2 18906 2669 18906 2669 0 net138
rlabel metal1 18078 2278 18078 2278 0 net139
rlabel metal1 36202 2414 36202 2414 0 net14
rlabel via2 18354 2907 18354 2907 0 net140
rlabel metal2 32430 2210 32430 2210 0 net141
rlabel metal2 19182 2227 19182 2227 0 net142
rlabel metal2 17342 1989 17342 1989 0 net143
rlabel metal2 33902 1700 33902 1700 0 net144
rlabel metal2 16698 1938 16698 1938 0 net145
rlabel metal1 2806 7378 2806 7378 0 net146
rlabel metal1 36938 2550 36938 2550 0 net15
rlabel metal4 36156 1836 36156 1836 0 net16
rlabel metal1 37812 2278 37812 2278 0 net17
rlabel metal2 38042 3910 38042 3910 0 net18
rlabel metal2 38318 2176 38318 2176 0 net19
rlabel metal1 38916 2278 38916 2278 0 net2
rlabel metal1 38594 1938 38594 1938 0 net20
rlabel metal2 5934 2312 5934 2312 0 net21
rlabel metal1 4922 1904 4922 1904 0 net22
rlabel metal1 5566 2040 5566 2040 0 net23
rlabel metal1 6302 2584 6302 2584 0 net24
rlabel metal1 8188 2278 8188 2278 0 net25
rlabel metal1 9430 2278 9430 2278 0 net26
rlabel metal2 9338 3366 9338 3366 0 net27
rlabel metal1 8786 2550 8786 2550 0 net28
rlabel metal1 9108 2550 9108 2550 0 net29
rlabel metal1 36754 2448 36754 2448 0 net3
rlabel metal2 9430 2023 9430 2023 0 net30
rlabel metal2 19458 2244 19458 2244 0 net31
rlabel metal2 9982 3264 9982 3264 0 net32
rlabel metal1 6164 2278 6164 2278 0 net33
rlabel metal2 6210 3570 6210 3570 0 net34
rlabel metal1 6578 1564 6578 1564 0 net35
rlabel metal2 6854 1836 6854 1836 0 net36
rlabel metal1 17066 2516 17066 2516 0 net37
rlabel metal1 21574 1802 21574 1802 0 net38
rlabel metal1 7682 2312 7682 2312 0 net39
rlabel metal1 37352 2890 37352 2890 0 net4
rlabel metal2 16974 2278 16974 2278 0 net40
rlabel metal2 10258 3638 10258 3638 0 net41
rlabel metal1 13248 2550 13248 2550 0 net42
rlabel metal1 13938 2278 13938 2278 0 net43
rlabel metal2 13938 3604 13938 3604 0 net44
rlabel metal1 19504 1870 19504 1870 0 net45
rlabel metal1 19550 2550 19550 2550 0 net46
rlabel metal2 15134 3264 15134 3264 0 net47
rlabel metal2 10534 1921 10534 1921 0 net48
rlabel metal2 10810 1717 10810 1717 0 net49
rlabel metal1 38502 1972 38502 1972 0 net5
rlabel metal2 11086 3111 11086 3111 0 net50
rlabel metal1 17986 1870 17986 1870 0 net51
rlabel metal2 13294 2227 13294 2227 0 net52
rlabel metal2 12006 3281 12006 3281 0 net53
rlabel metal3 18676 2448 18676 2448 0 net54
rlabel metal2 12558 3009 12558 3009 0 net55
rlabel metal2 12834 1972 12834 1972 0 net56
rlabel metal1 13754 2482 13754 2482 0 net57
rlabel metal1 17894 2958 17894 2958 0 net58
rlabel metal1 17710 2618 17710 2618 0 net59
rlabel metal1 40204 2550 40204 2550 0 net6
rlabel metal2 17802 2587 17802 2587 0 net60
rlabel metal1 18768 3026 18768 3026 0 net61
rlabel metal1 18998 2992 18998 2992 0 net62
rlabel metal1 19320 3026 19320 3026 0 net63
rlabel metal1 14996 2414 14996 2414 0 net64
rlabel metal1 15272 2414 15272 2414 0 net65
rlabel metal1 15548 2414 15548 2414 0 net66
rlabel metal1 15824 2414 15824 2414 0 net67
rlabel metal1 16100 2414 16100 2414 0 net68
rlabel metal1 16606 3366 16606 3366 0 net69
rlabel metal2 40158 2788 40158 2788 0 net7
rlabel metal1 17066 2992 17066 2992 0 net70
rlabel metal1 17066 3638 17066 3638 0 net71
rlabel metal1 17158 2414 17158 2414 0 net72
rlabel metal1 33948 2618 33948 2618 0 net73
rlabel metal1 17250 7412 17250 7412 0 net74
rlabel metal2 24886 6630 24886 6630 0 net75
rlabel metal1 27324 7446 27324 7446 0 net76
rlabel metal1 29118 3706 29118 3706 0 net77
rlabel metal2 31786 4998 31786 4998 0 net78
rlabel metal1 37950 7480 37950 7480 0 net79
rlabel metal1 39284 2414 39284 2414 0 net8
rlabel metal2 35558 3060 35558 3060 0 net80
rlabel metal1 39652 2618 39652 2618 0 net81
rlabel metal1 40342 2618 40342 2618 0 net82
rlabel metal1 41492 2618 41492 2618 0 net83
rlabel metal1 43010 2618 43010 2618 0 net84
rlabel metal2 5750 6800 5750 6800 0 net85
rlabel metal1 34822 3162 34822 3162 0 net86
rlabel metal2 35006 2006 35006 2006 0 net87
rlabel metal1 35512 3162 35512 3162 0 net88
rlabel metal1 14168 2618 14168 2618 0 net89
rlabel metal1 40526 2414 40526 2414 0 net9
rlabel metal1 16698 5882 16698 5882 0 net90
rlabel metal1 18676 7446 18676 7446 0 net91
rlabel metal1 20562 7480 20562 7480 0 net92
rlabel metal1 23184 6630 23184 6630 0 net93
rlabel metal1 18124 2346 18124 2346 0 net94
rlabel metal1 18446 2550 18446 2550 0 net95
rlabel metal1 19136 2278 19136 2278 0 net96
rlabel metal1 19688 2414 19688 2414 0 net97
rlabel metal1 22770 2448 22770 2448 0 net98
rlabel metal1 23138 3094 23138 3094 0 net99
<< properties >>
string FIXED_BBOX 0 0 45000 10000
<< end >>
