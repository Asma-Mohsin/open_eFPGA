module DSP (Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    VGND,
    VPWR,
    Tile_X0Y0_E1BEG,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2BEG,
    Tile_X0Y0_E2BEGb,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6BEG,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4BEG,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_NN4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_SS4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W1END,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W2END,
    Tile_X0Y0_W2MID,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_W6END,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y0_WW4END,
    Tile_X0Y1_E1BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2BEG,
    Tile_X0Y1_E2BEGb,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6BEG,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4BEG,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_NN4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_SS4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W1END,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W2END,
    Tile_X0Y1_W2MID,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_W6END,
    Tile_X0Y1_WW4BEG,
    Tile_X0Y1_WW4END);
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 input VGND;
 input VPWR;
 output [3:0] Tile_X0Y0_E1BEG;
 input [3:0] Tile_X0Y0_E1END;
 output [7:0] Tile_X0Y0_E2BEG;
 output [7:0] Tile_X0Y0_E2BEGb;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 output [11:0] Tile_X0Y0_E6BEG;
 input [11:0] Tile_X0Y0_E6END;
 output [15:0] Tile_X0Y0_EE4BEG;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 output [15:0] Tile_X0Y0_NN4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 input [15:0] Tile_X0Y0_SS4END;
 output [3:0] Tile_X0Y0_W1BEG;
 input [3:0] Tile_X0Y0_W1END;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 input [7:0] Tile_X0Y0_W2END;
 input [7:0] Tile_X0Y0_W2MID;
 output [11:0] Tile_X0Y0_W6BEG;
 input [11:0] Tile_X0Y0_W6END;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [15:0] Tile_X0Y0_WW4END;
 output [3:0] Tile_X0Y1_E1BEG;
 input [3:0] Tile_X0Y1_E1END;
 output [7:0] Tile_X0Y1_E2BEG;
 output [7:0] Tile_X0Y1_E2BEGb;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 output [11:0] Tile_X0Y1_E6BEG;
 input [11:0] Tile_X0Y1_E6END;
 output [15:0] Tile_X0Y1_EE4BEG;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 input [15:0] Tile_X0Y1_NN4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [15:0] Tile_X0Y1_SS4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 input [3:0] Tile_X0Y1_W1END;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 input [7:0] Tile_X0Y1_W2END;
 input [7:0] Tile_X0Y1_W2MID;
 output [11:0] Tile_X0Y1_W6BEG;
 input [11:0] Tile_X0Y1_W6END;
 output [15:0] Tile_X0Y1_WW4BEG;
 input [15:0] Tile_X0Y1_WW4END;

 wire \Tile_X0Y0_DSP_top/ConfigBits[0] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[100] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[101] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[102] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[103] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[104] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[105] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[106] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[107] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[108] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[109] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[10] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[110] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[111] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[112] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[113] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[114] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[115] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[116] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[117] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[118] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[119] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[11] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[120] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[121] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[122] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[123] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[124] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[125] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[126] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[127] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[128] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[129] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[12] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[130] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[131] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[132] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[133] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[134] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[135] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[136] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[137] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[138] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[139] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[13] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[140] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[141] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[142] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[143] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[144] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[145] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[146] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[147] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[148] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[149] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[14] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[150] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[151] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[152] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[153] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[154] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[155] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[156] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[157] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[158] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[159] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[15] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[160] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[161] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[162] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[163] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[164] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[165] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[166] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[167] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[168] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[169] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[16] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[170] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[171] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[172] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[173] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[174] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[175] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[176] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[177] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[178] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[179] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[17] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[180] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[181] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[182] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[183] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[184] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[185] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[186] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[187] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[188] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[189] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[18] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[190] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[191] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[192] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[193] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[194] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[195] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[196] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[197] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[198] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[199] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[19] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[1] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[200] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[201] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[202] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[203] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[204] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[205] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[206] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[207] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[208] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[209] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[20] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[210] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[211] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[212] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[213] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[214] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[215] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[216] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[217] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[218] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[219] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[21] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[220] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[221] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[222] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[223] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[224] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[225] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[226] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[227] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[228] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[229] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[22] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[230] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[231] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[232] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[233] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[234] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[235] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[236] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[237] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[238] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[239] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[23] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[240] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[241] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[242] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[243] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[244] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[245] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[246] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[247] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[248] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[249] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[24] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[250] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[251] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[252] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[253] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[254] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[255] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[256] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[257] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[258] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[259] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[25] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[260] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[261] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[262] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[263] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[264] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[265] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[266] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[267] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[268] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[269] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[26] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[270] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[271] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[272] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[273] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[274] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[275] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[276] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[277] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[278] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[279] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[27] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[280] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[281] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[282] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[283] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[284] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[285] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[286] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[287] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[288] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[289] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[28] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[290] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[291] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[292] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[293] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[294] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[295] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[296] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[297] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[298] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[299] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[29] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[2] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[300] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[301] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[302] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[303] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[304] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[305] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[306] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[307] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[308] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[309] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[30] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[310] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[311] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[312] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[313] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[314] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[315] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[316] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[317] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[318] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[319] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[31] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[320] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[321] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[322] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[323] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[324] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[325] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[326] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[327] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[328] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[329] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[32] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[330] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[331] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[332] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[333] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[334] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[335] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[336] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[337] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[338] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[339] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[33] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[340] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[341] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[342] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[343] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[344] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[345] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[346] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[347] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[348] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[349] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[34] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[350] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[351] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[352] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[353] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[354] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[355] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[356] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[357] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[358] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[359] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[35] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[360] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[361] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[362] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[363] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[364] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[365] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[366] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[367] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[368] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[369] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[36] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[370] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[371] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[372] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[373] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[374] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[375] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[376] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[377] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[378] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[379] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[37] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[380] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[381] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[382] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[383] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[384] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[385] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[386] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[387] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[388] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[389] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[38] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[390] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[391] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[392] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[393] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[394] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[395] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[396] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[397] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[398] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[399] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[39] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[3] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[400] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[401] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[402] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[403] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[404] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[405] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[40] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[41] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[42] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[43] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[44] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[45] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[46] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[47] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[48] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[49] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[4] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[50] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[51] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[52] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[53] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[54] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[55] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[56] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[57] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[58] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[59] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[5] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[60] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[61] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[62] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[63] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[64] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[65] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[66] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[67] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[68] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[69] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[6] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[70] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[71] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[72] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[73] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[74] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[75] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[76] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[77] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[78] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[79] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[7] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[80] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[81] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[82] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[83] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[84] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[85] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[86] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[87] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[88] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[89] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[8] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[90] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[91] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[92] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[93] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[94] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[95] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[96] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[97] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[98] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[99] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[9] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[0] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[100] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[101] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[102] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[103] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[104] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[105] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[106] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[107] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[108] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[109] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[10] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[110] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[111] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[112] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[113] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[114] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[115] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[116] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[117] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[118] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[119] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[11] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[120] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[121] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[122] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[123] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[124] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[125] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[126] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[127] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[128] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[129] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[12] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[130] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[131] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[132] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[133] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[134] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[135] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[136] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[137] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[138] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[139] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[13] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[140] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[141] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[142] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[143] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[144] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[145] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[146] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[147] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[148] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[149] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[14] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[150] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[151] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[152] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[153] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[154] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[155] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[156] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[157] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[158] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[159] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[15] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[160] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[161] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[162] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[163] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[164] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[165] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[166] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[167] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[168] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[169] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[16] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[170] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[171] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[172] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[173] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[174] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[175] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[176] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[177] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[178] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[179] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[17] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[180] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[181] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[182] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[183] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[184] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[185] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[186] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[187] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[188] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[189] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[18] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[190] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[191] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[192] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[193] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[194] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[195] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[196] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[197] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[198] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[199] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[19] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[1] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[200] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[201] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[202] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[203] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[204] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[205] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[206] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[207] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[208] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[209] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[20] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[210] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[211] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[212] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[213] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[214] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[215] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[216] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[217] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[218] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[219] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[21] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[220] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[221] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[222] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[223] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[224] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[225] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[226] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[227] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[228] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[229] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[22] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[230] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[231] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[232] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[233] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[234] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[235] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[236] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[237] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[238] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[239] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[23] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[240] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[241] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[242] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[243] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[244] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[245] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[246] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[247] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[248] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[249] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[24] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[250] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[251] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[252] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[253] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[254] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[255] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[256] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[257] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[258] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[259] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[25] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[260] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[261] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[262] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[263] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[264] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[265] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[266] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[267] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[268] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[269] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[26] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[270] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[271] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[272] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[273] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[274] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[275] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[276] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[277] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[278] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[279] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[27] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[280] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[281] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[282] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[283] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[284] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[285] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[286] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[287] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[288] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[289] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[28] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[290] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[291] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[292] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[293] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[294] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[295] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[296] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[297] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[298] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[299] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[29] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[2] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[300] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[301] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[302] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[303] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[304] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[305] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[306] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[307] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[308] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[309] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[30] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[310] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[311] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[312] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[313] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[314] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[315] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[316] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[317] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[318] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[319] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[31] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[320] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[321] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[322] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[323] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[324] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[325] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[326] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[327] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[328] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[329] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[32] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[330] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[331] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[332] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[333] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[334] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[335] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[336] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[337] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[338] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[339] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[33] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[340] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[341] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[342] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[343] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[344] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[345] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[346] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[347] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[348] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[349] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[34] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[350] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[351] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[352] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[353] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[354] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[355] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[356] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[357] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[358] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[359] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[35] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[360] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[361] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[362] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[363] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[364] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[365] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[366] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[367] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[368] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[369] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[36] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[370] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[371] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[372] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[373] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[374] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[375] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[376] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[377] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[378] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[379] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[37] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[380] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[381] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[382] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[383] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[384] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[385] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[386] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[387] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[388] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[389] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[38] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[390] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[391] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[392] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[393] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[394] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[395] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[396] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[397] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[398] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[399] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[39] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[3] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[400] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[401] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[402] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[403] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[404] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[405] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[40] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[41] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[42] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[43] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[44] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[45] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[46] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[47] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[48] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[49] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[4] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[50] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[51] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[52] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[53] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[54] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[55] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[56] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[57] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[58] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[59] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[5] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[60] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[61] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[62] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[63] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[64] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[65] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[66] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[67] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[68] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[69] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[6] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[70] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[71] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[72] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[73] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[74] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[75] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[76] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[77] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[78] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[79] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[7] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[80] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[81] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[82] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[83] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[84] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[85] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[86] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[87] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[88] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[89] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[8] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[90] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[91] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[92] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[93] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[94] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[95] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[96] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[97] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[98] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[99] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[9] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[0] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[10] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[11] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[12] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[13] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[14] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[15] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[16] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[17] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[18] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[19] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[1] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[20] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[21] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[22] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[23] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[24] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[25] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[26] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[27] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[28] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[29] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[2] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[30] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[31] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[3] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[4] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[5] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[6] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[7] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[8] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[9] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[0] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[10] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[11] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[12] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[13] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[14] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[15] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[16] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[17] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[18] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[19] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[1] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[2] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[3] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[4] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[5] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[6] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[7] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[8] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[9] ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/J2END_AB_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2END_AB_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2END_AB_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2END_AB_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2END_CD_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2END_CD_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2END_CD_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2END_CD_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2END_EF_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2END_EF_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2END_EF_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2END_EF_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2END_GH_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2END_GH_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2END_GH_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABa_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABa_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABa_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABb_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABb_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDa_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDa_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDa_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDb_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDb_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFa_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFa_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFa_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFb_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFb_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHa_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHa_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHa_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHb_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHb_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHb_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[0] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[1] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[2] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[4] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[5] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[6] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[7] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[0] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[1] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[2] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[4] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[5] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[6] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[7] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[0] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[1] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[2] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[4] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[5] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[6] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[7] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[0] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[1] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[2] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[4] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[5] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[6] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[7] ;
 wire \Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J_l_AB_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J_l_AB_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J_l_AB_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J_l_CD_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J_l_CD_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J_l_CD_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J_l_EF_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J_l_EF_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J_l_EF_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J_l_GH_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J_l_GH_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J_l_GH_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[9] ;
 wire \Tile_X0Y0_S1BEG[0] ;
 wire \Tile_X0Y0_S1BEG[1] ;
 wire \Tile_X0Y0_S1BEG[2] ;
 wire \Tile_X0Y0_S1BEG[3] ;
 wire \Tile_X0Y0_S2BEG[0] ;
 wire \Tile_X0Y0_S2BEG[1] ;
 wire \Tile_X0Y0_S2BEG[2] ;
 wire \Tile_X0Y0_S2BEG[3] ;
 wire \Tile_X0Y0_S2BEG[4] ;
 wire \Tile_X0Y0_S2BEG[5] ;
 wire \Tile_X0Y0_S2BEG[6] ;
 wire \Tile_X0Y0_S2BEG[7] ;
 wire \Tile_X0Y0_S2BEGb[0] ;
 wire \Tile_X0Y0_S2BEGb[1] ;
 wire \Tile_X0Y0_S2BEGb[2] ;
 wire \Tile_X0Y0_S2BEGb[3] ;
 wire \Tile_X0Y0_S2BEGb[4] ;
 wire \Tile_X0Y0_S2BEGb[5] ;
 wire \Tile_X0Y0_S2BEGb[6] ;
 wire \Tile_X0Y0_S2BEGb[7] ;
 wire \Tile_X0Y0_S4BEG[0] ;
 wire \Tile_X0Y0_S4BEG[10] ;
 wire \Tile_X0Y0_S4BEG[11] ;
 wire \Tile_X0Y0_S4BEG[12] ;
 wire \Tile_X0Y0_S4BEG[13] ;
 wire \Tile_X0Y0_S4BEG[14] ;
 wire \Tile_X0Y0_S4BEG[15] ;
 wire \Tile_X0Y0_S4BEG[1] ;
 wire \Tile_X0Y0_S4BEG[2] ;
 wire \Tile_X0Y0_S4BEG[3] ;
 wire \Tile_X0Y0_S4BEG[4] ;
 wire \Tile_X0Y0_S4BEG[5] ;
 wire \Tile_X0Y0_S4BEG[6] ;
 wire \Tile_X0Y0_S4BEG[7] ;
 wire \Tile_X0Y0_S4BEG[8] ;
 wire \Tile_X0Y0_S4BEG[9] ;
 wire \Tile_X0Y0_SS4BEG[0] ;
 wire \Tile_X0Y0_SS4BEG[10] ;
 wire \Tile_X0Y0_SS4BEG[11] ;
 wire \Tile_X0Y0_SS4BEG[12] ;
 wire \Tile_X0Y0_SS4BEG[13] ;
 wire \Tile_X0Y0_SS4BEG[14] ;
 wire \Tile_X0Y0_SS4BEG[15] ;
 wire \Tile_X0Y0_SS4BEG[1] ;
 wire \Tile_X0Y0_SS4BEG[2] ;
 wire \Tile_X0Y0_SS4BEG[3] ;
 wire \Tile_X0Y0_SS4BEG[4] ;
 wire \Tile_X0Y0_SS4BEG[5] ;
 wire \Tile_X0Y0_SS4BEG[6] ;
 wire \Tile_X0Y0_SS4BEG[7] ;
 wire \Tile_X0Y0_SS4BEG[8] ;
 wire \Tile_X0Y0_SS4BEG[9] ;
 wire \Tile_X0Y0_top2bot[0] ;
 wire \Tile_X0Y0_top2bot[10] ;
 wire \Tile_X0Y0_top2bot[11] ;
 wire \Tile_X0Y0_top2bot[12] ;
 wire \Tile_X0Y0_top2bot[13] ;
 wire \Tile_X0Y0_top2bot[14] ;
 wire \Tile_X0Y0_top2bot[15] ;
 wire \Tile_X0Y0_top2bot[16] ;
 wire \Tile_X0Y0_top2bot[17] ;
 wire \Tile_X0Y0_top2bot[1] ;
 wire \Tile_X0Y0_top2bot[2] ;
 wire \Tile_X0Y0_top2bot[3] ;
 wire \Tile_X0Y0_top2bot[4] ;
 wire \Tile_X0Y0_top2bot[5] ;
 wire \Tile_X0Y0_top2bot[6] ;
 wire \Tile_X0Y0_top2bot[7] ;
 wire \Tile_X0Y0_top2bot[8] ;
 wire \Tile_X0Y0_top2bot[9] ;
 wire \Tile_X0Y1_DSP_bot/A0 ;
 wire \Tile_X0Y1_DSP_bot/A1 ;
 wire \Tile_X0Y1_DSP_bot/A2 ;
 wire \Tile_X0Y1_DSP_bot/A3 ;
 wire \Tile_X0Y1_DSP_bot/A4 ;
 wire \Tile_X0Y1_DSP_bot/A5 ;
 wire \Tile_X0Y1_DSP_bot/A6 ;
 wire \Tile_X0Y1_DSP_bot/A7 ;
 wire \Tile_X0Y1_DSP_bot/B0 ;
 wire \Tile_X0Y1_DSP_bot/B1 ;
 wire \Tile_X0Y1_DSP_bot/B2 ;
 wire \Tile_X0Y1_DSP_bot/B3 ;
 wire \Tile_X0Y1_DSP_bot/B4 ;
 wire \Tile_X0Y1_DSP_bot/B5 ;
 wire \Tile_X0Y1_DSP_bot/B6 ;
 wire \Tile_X0Y1_DSP_bot/B7 ;
 wire \Tile_X0Y1_DSP_bot/C0 ;
 wire \Tile_X0Y1_DSP_bot/C1 ;
 wire \Tile_X0Y1_DSP_bot/C10 ;
 wire \Tile_X0Y1_DSP_bot/C11 ;
 wire \Tile_X0Y1_DSP_bot/C12 ;
 wire \Tile_X0Y1_DSP_bot/C13 ;
 wire \Tile_X0Y1_DSP_bot/C14 ;
 wire \Tile_X0Y1_DSP_bot/C15 ;
 wire \Tile_X0Y1_DSP_bot/C16 ;
 wire \Tile_X0Y1_DSP_bot/C17 ;
 wire \Tile_X0Y1_DSP_bot/C18 ;
 wire \Tile_X0Y1_DSP_bot/C19 ;
 wire \Tile_X0Y1_DSP_bot/C2 ;
 wire \Tile_X0Y1_DSP_bot/C3 ;
 wire \Tile_X0Y1_DSP_bot/C4 ;
 wire \Tile_X0Y1_DSP_bot/C5 ;
 wire \Tile_X0Y1_DSP_bot/C6 ;
 wire \Tile_X0Y1_DSP_bot/C7 ;
 wire \Tile_X0Y1_DSP_bot/C8 ;
 wire \Tile_X0Y1_DSP_bot/C9 ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[0] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[100] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[101] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[102] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[103] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[104] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[105] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[106] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[107] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[108] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[109] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[10] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[110] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[111] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[112] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[113] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[114] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[115] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[116] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[117] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[118] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[119] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[11] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[120] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[121] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[122] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[123] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[124] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[125] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[126] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[127] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[128] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[129] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[12] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[130] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[131] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[132] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[133] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[134] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[135] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[136] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[137] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[138] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[139] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[13] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[140] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[141] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[142] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[143] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[144] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[145] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[146] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[147] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[148] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[149] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[14] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[150] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[151] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[152] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[153] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[154] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[155] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[156] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[157] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[158] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[159] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[15] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[160] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[161] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[162] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[163] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[164] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[165] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[166] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[167] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[168] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[169] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[16] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[170] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[171] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[172] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[173] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[174] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[175] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[176] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[177] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[178] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[179] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[17] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[180] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[181] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[182] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[183] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[184] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[185] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[186] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[187] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[188] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[189] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[18] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[190] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[191] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[192] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[193] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[194] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[195] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[196] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[197] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[198] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[199] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[19] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[1] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[200] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[201] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[202] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[203] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[204] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[205] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[206] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[207] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[208] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[209] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[20] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[210] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[211] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[212] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[213] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[214] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[215] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[216] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[217] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[218] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[219] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[21] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[220] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[221] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[222] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[223] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[224] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[225] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[226] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[227] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[228] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[229] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[22] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[230] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[231] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[232] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[233] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[234] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[235] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[236] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[237] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[238] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[239] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[23] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[240] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[241] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[242] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[243] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[244] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[245] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[246] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[247] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[248] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[249] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[24] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[250] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[251] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[252] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[253] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[254] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[255] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[256] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[257] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[258] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[259] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[25] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[260] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[261] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[262] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[263] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[264] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[265] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[266] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[267] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[268] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[269] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[26] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[270] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[271] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[272] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[273] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[274] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[275] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[276] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[277] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[278] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[279] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[27] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[280] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[281] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[282] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[283] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[284] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[285] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[286] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[287] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[288] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[289] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[28] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[290] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[291] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[292] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[293] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[294] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[295] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[296] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[297] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[298] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[299] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[29] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[2] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[300] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[301] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[302] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[303] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[304] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[305] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[306] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[307] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[308] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[309] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[30] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[310] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[311] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[312] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[313] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[314] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[315] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[316] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[317] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[318] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[319] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[31] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[320] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[321] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[322] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[323] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[324] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[325] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[326] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[327] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[328] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[329] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[32] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[330] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[331] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[332] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[333] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[334] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[335] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[336] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[337] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[338] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[339] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[33] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[340] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[341] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[342] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[343] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[344] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[345] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[346] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[347] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[348] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[349] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[34] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[350] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[351] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[352] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[353] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[354] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[355] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[356] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[357] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[358] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[359] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[35] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[360] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[361] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[362] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[363] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[364] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[365] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[366] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[367] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[368] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[369] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[36] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[370] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[371] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[372] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[373] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[374] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[375] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[376] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[377] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[378] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[379] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[37] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[380] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[381] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[382] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[383] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[384] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[385] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[386] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[387] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[388] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[389] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[38] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[390] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[391] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[392] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[393] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[394] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[395] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[396] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[397] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[398] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[399] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[39] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[3] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[400] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[401] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[402] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[403] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[404] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[405] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[406] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[407] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[408] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[409] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[40] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[410] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[411] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[412] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[413] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[414] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[415] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[41] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[42] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[43] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[44] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[45] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[46] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[47] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[48] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[49] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[4] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[50] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[51] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[52] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[53] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[54] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[55] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[56] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[57] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[58] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[59] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[5] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[60] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[61] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[62] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[63] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[64] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[65] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[66] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[67] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[68] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[69] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[6] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[70] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[71] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[72] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[73] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[74] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[75] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[76] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[77] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[78] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[79] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[7] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[80] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[81] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[82] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[83] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[84] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[85] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[86] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[87] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[88] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[89] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[8] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[90] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[91] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[92] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[93] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[94] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[95] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[96] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[97] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[98] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[99] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[9] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[0] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[100] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[101] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[102] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[103] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[104] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[105] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[106] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[107] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[108] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[109] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[10] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[110] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[111] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[112] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[113] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[114] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[115] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[116] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[117] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[118] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[119] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[11] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[120] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[121] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[122] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[123] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[124] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[125] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[126] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[127] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[128] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[129] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[12] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[130] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[131] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[132] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[133] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[134] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[135] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[136] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[137] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[138] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[139] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[13] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[140] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[141] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[142] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[143] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[144] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[145] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[146] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[147] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[148] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[149] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[14] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[150] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[151] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[152] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[153] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[154] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[155] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[156] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[157] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[158] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[159] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[15] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[160] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[161] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[162] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[163] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[164] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[165] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[166] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[167] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[168] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[169] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[16] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[170] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[171] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[172] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[173] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[174] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[175] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[176] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[177] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[178] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[179] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[17] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[180] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[181] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[182] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[183] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[184] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[185] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[186] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[187] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[188] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[189] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[18] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[190] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[191] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[192] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[193] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[194] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[195] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[196] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[197] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[198] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[199] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[19] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[1] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[200] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[201] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[202] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[203] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[204] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[205] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[206] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[207] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[208] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[209] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[20] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[210] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[211] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[212] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[213] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[214] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[215] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[216] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[217] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[218] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[219] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[21] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[220] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[221] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[222] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[223] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[224] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[225] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[226] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[227] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[228] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[229] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[22] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[230] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[231] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[232] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[233] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[234] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[235] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[236] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[237] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[238] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[239] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[23] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[240] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[241] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[242] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[243] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[244] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[245] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[246] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[247] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[248] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[249] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[24] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[250] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[251] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[252] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[253] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[254] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[255] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[256] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[257] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[258] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[259] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[25] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[260] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[261] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[262] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[263] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[264] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[265] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[266] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[267] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[268] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[269] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[26] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[270] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[271] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[272] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[273] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[274] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[275] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[276] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[277] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[278] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[279] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[27] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[280] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[281] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[282] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[283] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[284] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[285] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[286] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[287] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[288] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[289] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[28] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[290] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[291] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[292] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[293] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[294] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[295] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[296] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[297] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[298] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[299] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[29] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[2] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[300] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[301] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[302] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[303] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[304] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[305] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[306] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[307] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[308] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[309] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[30] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[310] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[311] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[312] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[313] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[314] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[315] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[316] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[317] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[318] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[319] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[31] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[320] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[321] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[322] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[323] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[324] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[325] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[326] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[327] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[328] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[329] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[32] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[330] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[331] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[332] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[333] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[334] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[335] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[336] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[337] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[338] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[339] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[33] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[340] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[341] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[342] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[343] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[344] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[345] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[346] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[347] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[348] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[349] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[34] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[350] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[351] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[352] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[353] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[354] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[355] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[356] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[357] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[358] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[359] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[35] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[360] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[361] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[362] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[363] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[364] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[365] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[366] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[367] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[368] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[369] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[36] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[370] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[371] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[372] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[373] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[374] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[375] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[376] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[377] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[378] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[379] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[37] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[380] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[381] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[382] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[383] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[384] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[385] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[386] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[387] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[388] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[389] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[38] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[390] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[391] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[392] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[393] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[394] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[395] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[396] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[397] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[398] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[399] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[39] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[3] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[400] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[401] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[402] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[403] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[404] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[405] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[406] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[407] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[408] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[409] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[40] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[410] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[411] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[412] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[413] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[414] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[415] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[41] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[42] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[43] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[44] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[45] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[46] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[47] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[48] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[49] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[4] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[50] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[51] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[52] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[53] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[54] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[55] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[56] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[57] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[58] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[59] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[5] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[60] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[61] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[62] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[63] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[64] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[65] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[66] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[67] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[68] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[69] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[6] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[70] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[71] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[72] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[73] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[74] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[75] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[76] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[77] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[78] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[79] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[7] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[80] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[81] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[82] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[83] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[84] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[85] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[86] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[87] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[88] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[89] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[8] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[90] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[91] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[92] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[93] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[94] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[95] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[96] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[97] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[98] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[99] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[9] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[0] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[10] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[11] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[12] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[13] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[14] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[15] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[16] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[17] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[18] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[19] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[1] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[20] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[21] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[22] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[23] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[24] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[25] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[26] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[27] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[28] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[29] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[2] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[30] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[31] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[3] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[4] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[5] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[6] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[7] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[8] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[9] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[0] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[10] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[11] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[12] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[13] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[14] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[15] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[16] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[17] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[18] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[19] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[1] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[2] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[3] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[4] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[5] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[6] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[7] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[8] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[9] ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[0] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[10] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[11] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[12] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[13] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[14] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[15] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[16] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[18] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[19] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[1] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[2] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[3] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[4] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[5] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[6] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[7] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[8] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[9] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[0] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[1] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[2] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[5] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[6] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[7] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[0] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[1] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[3] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[4] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[5] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[6] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[7] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[0] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[10] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[11] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[12] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[13] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[14] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[15] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[16] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[17] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[18] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[19] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[1] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[2] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[3] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[4] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[5] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[6] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[7] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[8] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[9] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0000_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0001_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0002_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0003_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0004_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0005_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0006_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0007_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0008_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0009_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0010_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0011_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0012_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0013_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0014_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0015_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0016_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0017_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0018_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0019_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0020_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0022_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0023_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0031_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0035_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0036_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0039_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0042_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0043_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0053_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0055_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0056_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0057_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0058_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0059_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0060_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0061_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0062_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0066_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0068_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0069_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0072_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0077_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0078_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0081_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0083_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0084_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0087_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0088_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0089_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0090_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0091_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0092_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0093_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0095_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0096_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0097_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0098_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0099_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0100_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0104_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0110_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0111_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0115_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0116_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0118_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0119_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0120_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0126_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0128_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0129_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0130_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0131_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0133_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0134_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0139_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0140_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0144_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0148_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0150_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0153_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0156_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0160_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0161_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0162_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0167_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0168_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0169_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0170_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0172_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0173_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0174_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0175_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0177_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0179_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0180_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0181_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0182_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0183_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0186_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0187_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0200_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0201_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0202_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0203_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0209_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0210_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0211_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0212_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0218_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0219_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0220_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0224_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0225_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0229_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0232_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0233_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0234_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0236_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0237_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0240_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0241_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0242_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0243_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0244_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0245_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0246_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0247_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0248_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0249_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0251_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0252_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0253_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0254_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0256_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0257_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0260_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0262_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0264_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0266_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0276_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0277_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0278_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0279_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0280_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0281_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0287_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0288_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0296_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0302_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0308_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0310_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0311_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0312_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0314_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0315_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0316_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0317_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0320_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0322_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0323_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0324_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0326_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0328_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0329_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0330_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0332_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0333_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0334_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0335_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0336_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0337_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0338_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0339_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0340_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0344_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0350_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0352_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0354_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0355_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0356_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0361_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0362_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0363_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0364_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0367_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0373_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0374_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0376_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0384_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0385_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0386_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0388_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0392_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0393_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0394_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0399_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0400_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0401_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0402_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0403_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0404_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0405_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0406_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0408_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0412_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0413_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0418_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0419_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0420_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0421_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0422_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0425_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0426_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0427_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0429_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0430_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0431_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0432_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0433_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0434_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0436_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0437_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0441_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0447_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0456_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0458_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0459_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0462_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0465_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0468_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0469_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0470_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0471_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0474_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0475_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0477_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0479_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0480_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0481_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0482_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0485_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0486_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0487_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0489_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0495_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0499_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0500_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0502_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0503_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0504_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0505_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0506_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0507_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0508_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0509_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0510_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0511_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0512_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0513_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0514_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0515_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0517_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0518_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0520_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0522_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0524_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0526_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0528_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0530_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0531_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0532_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0537_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0538_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0540_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0541_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0542_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0544_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0546_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0547_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0548_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0550_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0551_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0553_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0555_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0556_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0558_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0559_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0565_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0566_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0567_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0568_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0571_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0572_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0574_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0575_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0576_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0577_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0578_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0580_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0582_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0583_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0584_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0585_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0587_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0588_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0589_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0590_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0592_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0593_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0595_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0600_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0601_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0602_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0605_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0606_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0608_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0615_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0616_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0617_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0618_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0619_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0620_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0621_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0622_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0627_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0628_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0629_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0630_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0631_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0633_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0635_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0636_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0637_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0638_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0640_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0642_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0643_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0644_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0645_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0647_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0648_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0649_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0650_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0651_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0652_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0653_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0654_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0655_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0659_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0661_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0662_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0665_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0666_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0668_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0674_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0675_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0676_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0678_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0680_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0684_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0685_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0686_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0687_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0688_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0689_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0690_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0691_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0693_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0694_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0698_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0700_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0703_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0704_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0705_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0706_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0708_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0709_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0710_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0712_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0715_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0716_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0717_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0718_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0719_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0720_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0721_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0722_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0723_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0724_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0726_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0727_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0729_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0731_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0732_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0735_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0736_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0737_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0738_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0739_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0740_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0742_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0743_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0744_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0745_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0746_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0747_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0748_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0749_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0750_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0751_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0752_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0753_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0754_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0756_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0757_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0758_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0759_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0761_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0766_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0767_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0768_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0769_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0770_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0772_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0773_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0774_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0776_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0779_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0781_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0782_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0783_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0784_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0785_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0786_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0788_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0789_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0791_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0792_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0793_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0794_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0796_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0797_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0800_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0801_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0803_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0804_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0805_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0806_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0807_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0808_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0811_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0812_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0816_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0817_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0818_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0819_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0820_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0821_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0822_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0823_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0824_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0825_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0826_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0827_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0828_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0831_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0832_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0833_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0834_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0835_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0836_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0837_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0838_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0839_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0840_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0841_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0842_ ;
 wire \Tile_X0Y1_DSP_bot/J2END_AB_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2END_AB_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2END_AB_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2END_CD_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2END_CD_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2END_CD_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2END_CD_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2END_EF_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2END_EF_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2END_EF_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2END_GH_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2END_GH_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2END_GH_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2END_GH_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[4] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[5] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[6] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[7] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[4] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[5] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[6] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[7] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[4] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[5] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[6] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[7] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[4] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[5] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[6] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[7] ;
 wire \Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J_l_AB_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J_l_AB_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J_l_AB_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J_l_CD_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J_l_CD_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J_l_CD_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J_l_EF_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J_l_EF_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J_l_EF_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J_l_GH_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J_l_GH_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J_l_GH_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/Q0 ;
 wire \Tile_X0Y1_DSP_bot/Q1 ;
 wire \Tile_X0Y1_DSP_bot/Q10 ;
 wire \Tile_X0Y1_DSP_bot/Q11 ;
 wire \Tile_X0Y1_DSP_bot/Q12 ;
 wire \Tile_X0Y1_DSP_bot/Q13 ;
 wire \Tile_X0Y1_DSP_bot/Q14 ;
 wire \Tile_X0Y1_DSP_bot/Q15 ;
 wire \Tile_X0Y1_DSP_bot/Q16 ;
 wire \Tile_X0Y1_DSP_bot/Q17 ;
 wire \Tile_X0Y1_DSP_bot/Q18 ;
 wire \Tile_X0Y1_DSP_bot/Q19 ;
 wire \Tile_X0Y1_DSP_bot/Q2 ;
 wire \Tile_X0Y1_DSP_bot/Q3 ;
 wire \Tile_X0Y1_DSP_bot/Q4 ;
 wire \Tile_X0Y1_DSP_bot/Q5 ;
 wire \Tile_X0Y1_DSP_bot/Q6 ;
 wire \Tile_X0Y1_DSP_bot/Q7 ;
 wire \Tile_X0Y1_DSP_bot/Q8 ;
 wire \Tile_X0Y1_DSP_bot/Q9 ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/clr ;
 wire \Tile_X0Y1_FrameStrobe_O[0] ;
 wire \Tile_X0Y1_FrameStrobe_O[10] ;
 wire \Tile_X0Y1_FrameStrobe_O[11] ;
 wire \Tile_X0Y1_FrameStrobe_O[12] ;
 wire \Tile_X0Y1_FrameStrobe_O[13] ;
 wire \Tile_X0Y1_FrameStrobe_O[14] ;
 wire \Tile_X0Y1_FrameStrobe_O[15] ;
 wire \Tile_X0Y1_FrameStrobe_O[16] ;
 wire \Tile_X0Y1_FrameStrobe_O[17] ;
 wire \Tile_X0Y1_FrameStrobe_O[18] ;
 wire \Tile_X0Y1_FrameStrobe_O[19] ;
 wire \Tile_X0Y1_FrameStrobe_O[1] ;
 wire \Tile_X0Y1_FrameStrobe_O[2] ;
 wire \Tile_X0Y1_FrameStrobe_O[3] ;
 wire \Tile_X0Y1_FrameStrobe_O[4] ;
 wire \Tile_X0Y1_FrameStrobe_O[5] ;
 wire \Tile_X0Y1_FrameStrobe_O[6] ;
 wire \Tile_X0Y1_FrameStrobe_O[7] ;
 wire \Tile_X0Y1_FrameStrobe_O[8] ;
 wire \Tile_X0Y1_FrameStrobe_O[9] ;
 wire \Tile_X0Y1_N1BEG[0] ;
 wire \Tile_X0Y1_N1BEG[1] ;
 wire \Tile_X0Y1_N1BEG[2] ;
 wire \Tile_X0Y1_N1BEG[3] ;
 wire \Tile_X0Y1_N2BEG[0] ;
 wire \Tile_X0Y1_N2BEG[1] ;
 wire \Tile_X0Y1_N2BEG[2] ;
 wire \Tile_X0Y1_N2BEG[3] ;
 wire \Tile_X0Y1_N2BEG[4] ;
 wire \Tile_X0Y1_N2BEG[5] ;
 wire \Tile_X0Y1_N2BEG[6] ;
 wire \Tile_X0Y1_N2BEG[7] ;
 wire \Tile_X0Y1_N2BEGb[0] ;
 wire \Tile_X0Y1_N2BEGb[1] ;
 wire \Tile_X0Y1_N2BEGb[2] ;
 wire \Tile_X0Y1_N2BEGb[3] ;
 wire \Tile_X0Y1_N2BEGb[4] ;
 wire \Tile_X0Y1_N2BEGb[5] ;
 wire \Tile_X0Y1_N2BEGb[6] ;
 wire \Tile_X0Y1_N2BEGb[7] ;
 wire \Tile_X0Y1_N4BEG[0] ;
 wire \Tile_X0Y1_N4BEG[10] ;
 wire \Tile_X0Y1_N4BEG[11] ;
 wire \Tile_X0Y1_N4BEG[12] ;
 wire \Tile_X0Y1_N4BEG[13] ;
 wire \Tile_X0Y1_N4BEG[14] ;
 wire \Tile_X0Y1_N4BEG[15] ;
 wire \Tile_X0Y1_N4BEG[1] ;
 wire \Tile_X0Y1_N4BEG[2] ;
 wire \Tile_X0Y1_N4BEG[3] ;
 wire \Tile_X0Y1_N4BEG[4] ;
 wire \Tile_X0Y1_N4BEG[5] ;
 wire \Tile_X0Y1_N4BEG[6] ;
 wire \Tile_X0Y1_N4BEG[7] ;
 wire \Tile_X0Y1_N4BEG[8] ;
 wire \Tile_X0Y1_N4BEG[9] ;
 wire \Tile_X0Y1_NN4BEG[0] ;
 wire \Tile_X0Y1_NN4BEG[10] ;
 wire \Tile_X0Y1_NN4BEG[11] ;
 wire \Tile_X0Y1_NN4BEG[12] ;
 wire \Tile_X0Y1_NN4BEG[13] ;
 wire \Tile_X0Y1_NN4BEG[14] ;
 wire \Tile_X0Y1_NN4BEG[15] ;
 wire \Tile_X0Y1_NN4BEG[1] ;
 wire \Tile_X0Y1_NN4BEG[2] ;
 wire \Tile_X0Y1_NN4BEG[3] ;
 wire \Tile_X0Y1_NN4BEG[4] ;
 wire \Tile_X0Y1_NN4BEG[5] ;
 wire \Tile_X0Y1_NN4BEG[6] ;
 wire \Tile_X0Y1_NN4BEG[7] ;
 wire \Tile_X0Y1_NN4BEG[8] ;
 wire \Tile_X0Y1_NN4BEG[9] ;
 wire Tile_X0Y1_UserCLKo;
 wire \Tile_X0Y1_bot2top[0] ;
 wire \Tile_X0Y1_bot2top[1] ;
 wire \Tile_X0Y1_bot2top[2] ;
 wire \Tile_X0Y1_bot2top[3] ;
 wire \Tile_X0Y1_bot2top[4] ;
 wire \Tile_X0Y1_bot2top[5] ;
 wire \Tile_X0Y1_bot2top[6] ;
 wire \Tile_X0Y1_bot2top[7] ;
 wire \Tile_X0Y1_bot2top[8] ;
 wire \Tile_X0Y1_bot2top[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\Tile_X0Y0_S2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\Tile_X0Y0_SS4BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(\Tile_X0Y1_DSP_bot/N4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(\Tile_X0Y1_DSP_bot/NN4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\Tile_X0Y0_SS4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\Tile_X0Y0_SS4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net283),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net295),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net341),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net345),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\Tile_X0Y0_SS4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net482),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net703),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net715),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(\Tile_X0Y0_SS4BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(\Tile_X0Y0_SS4BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\Tile_X0Y0_SS4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(\Tile_X0Y1_N1BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(\Tile_X0Y1_N1BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(\Tile_X0Y1_N1BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\Tile_X0Y0_SS4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(\Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(\Tile_X0Y0_DSP_top/JW2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(\Tile_X0Y1_DSP_bot/EE4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\Tile_X0Y0_SS4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(\Tile_X0Y1_DSP_bot/N4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\Tile_X0Y0_SS4BEG[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net665),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(\Tile_X0Y0_S1BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(\Tile_X0Y1_N1BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(\Tile_X0Y1_N1BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(\Tile_X0Y1_N1BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\Tile_X0Y0_SS4BEG[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\Tile_X0Y0_SS4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\Tile_X0Y0_SS4BEG[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\Tile_X0Y0_SS4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\Tile_X0Y0_SS4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\Tile_X0Y0_SS4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\Tile_X0Y0_SS4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\Tile_X0Y0_SS4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\Tile_X0Y1_FrameStrobe_O[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\Tile_X0Y1_FrameStrobe_O[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\Tile_X0Y1_FrameStrobe_O[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\Tile_X0Y1_FrameStrobe_O[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\Tile_X0Y1_FrameStrobe_O[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\Tile_X0Y0_SS4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\Tile_X0Y1_FrameStrobe_O[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\Tile_X0Y1_FrameStrobe_O[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\Tile_X0Y0_SS4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\Tile_X0Y1_FrameStrobe_O[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\Tile_X0Y1_FrameStrobe_O[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\Tile_X0Y1_FrameStrobe_O[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\Tile_X0Y1_FrameStrobe_O[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\Tile_X0Y1_FrameStrobe_O[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\Tile_X0Y1_FrameStrobe_O[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\Tile_X0Y1_FrameStrobe_O[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\Tile_X0Y1_FrameStrobe_O[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\Tile_X0Y1_FrameStrobe_O[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\Tile_X0Y1_FrameStrobe_O[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\Tile_X0Y0_SS4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\Tile_X0Y1_FrameStrobe_O[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\Tile_X0Y1_N1BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\Tile_X0Y1_N1BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\Tile_X0Y1_N1BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\Tile_X0Y1_N1BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\Tile_X0Y1_N1BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\Tile_X0Y1_N1BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\Tile_X0Y1_N1BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\Tile_X0Y1_N2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\Tile_X0Y0_DSP_top/E6BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\Tile_X0Y0_SS4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\Tile_X0Y0_DSP_top/EE4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\Tile_X0Y0_DSP_top/EE4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\Tile_X0Y0_DSP_top/JN2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\Tile_X0Y0_SS4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\Tile_X0Y0_SS4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\Tile_X0Y0_DSP_top/W6BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\Tile_X0Y0_SS4BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(\Tile_X0Y0_DSP_top/WW4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(\Tile_X0Y1_DSP_bot/B2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(\Tile_X0Y1_DSP_bot/E6BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(\Tile_X0Y1_DSP_bot/E6BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(\Tile_X0Y1_DSP_bot/E6BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(\Tile_X0Y1_DSP_bot/EE4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(\Tile_X0Y1_DSP_bot/EE4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(\Tile_X0Y1_DSP_bot/JE2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(\Tile_X0Y1_DSP_bot/JN2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(\Tile_X0Y1_DSP_bot/N4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_100_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_100_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_100_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_100_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_100_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_100_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_100_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_100_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_100_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_100_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_100_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_451 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_100_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_100_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_101_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_101_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_101_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_101_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_101_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_101_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_101_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_101_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_101_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_101_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_101_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_101_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_102_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_102_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_102_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_102_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_102_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_102_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_102_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_102_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_102_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_102_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_102_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_102_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_102_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_102_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_102_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_103_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_103_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_103_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_103_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_103_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_103_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_103_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_103_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_103_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_103_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_103_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_103_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_103_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_103_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_104_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_104_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_104_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_104_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_104_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_104_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_104_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_104_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_104_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_104_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_104_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_104_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_105_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_105_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_105_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_105_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_105_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_105_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_105_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_105_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_105_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_105_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_105_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_105_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_105_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_105_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_106_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_106_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_106_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_106_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_106_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_106_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_106_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_106_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_106_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_106_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_106_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_107_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_107_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_107_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_107_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_107_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_107_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_107_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_107_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_107_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_107_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_107_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_107_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_108_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_108_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_108_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_108_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_108_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_108_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_108_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_108_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_108_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_109_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_109_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_109_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_109_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_109_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_109_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_109_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_109_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_109_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_451 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_110_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_110_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_110_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_110_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_110_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_110_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_110_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_110_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_110_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_110_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_110_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_110_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_110_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_110_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_110_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_111_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_111_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_111_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_111_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_111_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_111_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_111_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_111_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_111_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_111_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_111_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_111_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_111_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_112_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_112_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_112_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_112_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_112_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_112_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_112_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_112_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_112_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_112_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_112_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_113_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_113_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_114_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_114_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_114_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_114_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_114_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_115_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_115_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_115_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_115_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_115_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_115_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_115_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_115_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_115_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_115_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_115_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_115_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_116_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_116_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_116_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_116_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_116_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_116_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_117_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_117_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_117_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_117_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_117_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_117_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_117_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_117_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_117_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_117_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_117_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_117_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_117_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_117_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_117_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_117_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_117_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_118_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_118_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_118_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_118_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_118_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_118_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_118_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_118_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_118_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_118_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_118_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_118_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_118_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_118_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_118_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_118_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_118_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_118_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_119_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_119_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_119_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_119_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_119_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_119_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_119_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_119_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_119_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_119_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_120_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_120_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_120_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_120_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_120_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_120_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_120_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_120_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_120_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_120_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_120_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_120_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_120_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_121_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_121_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_121_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_121_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_121_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_121_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_121_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_121_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_121_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_121_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_121_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_121_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_121_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_121_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_121_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_121_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_121_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_121_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_121_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_121_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_122_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_122_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_122_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_122_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_122_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_122_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_122_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_122_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_122_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_122_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_122_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_122_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_122_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_122_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_122_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_122_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_122_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_122_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_122_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_122_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_122_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_123_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_123_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_123_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_123_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_123_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_123_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_123_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_123_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_123_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_123_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_123_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_123_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_123_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_123_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_123_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_123_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_123_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_123_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_124_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_124_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_124_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_124_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_124_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_124_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_124_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_124_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_124_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_124_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_124_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_124_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_124_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_124_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_124_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_124_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_124_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_124_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_124_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_125_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_125_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_125_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_125_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_125_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_125_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_125_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_125_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_125_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_125_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_125_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_125_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_125_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_125_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_125_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_125_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_125_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_125_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_125_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_125_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_125_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_125_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_125_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_126_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_126_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_126_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_126_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_126_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_126_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_126_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_126_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_126_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_126_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_126_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_126_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_126_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_126_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_126_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_127_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_127_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_127_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_127_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_127_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_127_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_127_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_127_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_127_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_127_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_127_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_127_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_127_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_127_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_127_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_127_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_127_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_127_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_127_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_128_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_128_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_128_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_128_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_128_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_128_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_128_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_128_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_128_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_128_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_129_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_129_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_129_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_129_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_129_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_129_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_129_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_129_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_129_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_129_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_129_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_129_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_129_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_129_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_129_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_129_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_129_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_129_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_129_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_129_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_129_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_129_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_129_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_129_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_129_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_129_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_129_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_129_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_129_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_129_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_129_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_130_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_130_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_130_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_130_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_130_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_130_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_130_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_130_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_130_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_130_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_130_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_130_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_130_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_130_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_130_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_130_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_130_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_130_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_130_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_130_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_131_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_131_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_131_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_131_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_131_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_131_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_131_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_131_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_131_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_131_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_131_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_131_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_131_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_131_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_131_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_131_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_131_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_131_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_131_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_131_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_131_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_131_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_132_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_132_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_132_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_132_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_132_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_132_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_132_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_132_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_132_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_132_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_132_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_132_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_132_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_132_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_132_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_132_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_132_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_132_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_132_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_133_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_133_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_133_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_133_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_133_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_133_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_133_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_133_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_133_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_133_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_133_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_133_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_133_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_133_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_133_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_133_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_133_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_133_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_133_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_133_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_134_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_134_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_134_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_134_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_134_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_134_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_134_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_134_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_134_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_134_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_134_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_134_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_134_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_134_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_134_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_135_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_135_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_135_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_135_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_135_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_135_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_135_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_135_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_135_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_135_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_135_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_135_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_135_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_135_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_136_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_136_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_136_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_136_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_136_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_136_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_136_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_136_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_136_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_136_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_136_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_136_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_136_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_136_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_137_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_137_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_137_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_137_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_137_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_137_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_137_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_137_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_137_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_137_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_137_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_137_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_137_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_137_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_137_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_138_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_138_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_138_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_138_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_138_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_138_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_138_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_138_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_138_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_138_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_138_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_138_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_138_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_138_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_138_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_138_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_138_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_138_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_139_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_139_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_139_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_139_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_139_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_139_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_139_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_139_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_139_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_139_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_139_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_139_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_139_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_139_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_139_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_139_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_139_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_139_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_139_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_140_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_140_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_140_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_140_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_140_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_140_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_140_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_140_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_140_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_140_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_140_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_140_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_140_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_140_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_140_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_140_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_140_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_140_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_140_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_140_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_140_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_140_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_140_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_140_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_141_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_141_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_141_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_141_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_141_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_141_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_141_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_141_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_141_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_141_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_141_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_141_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_141_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_142_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_142_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_142_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_142_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_142_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_142_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_142_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_142_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_142_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_142_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_142_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_142_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_142_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_142_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_142_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_142_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_143_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_143_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_143_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_143_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_143_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_143_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_143_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_143_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_143_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_143_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_143_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_143_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_143_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_143_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_143_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_143_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_143_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_144_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_144_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_144_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_144_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_144_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_144_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_144_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_144_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_144_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_144_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_144_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_144_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_144_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_144_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_144_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_145_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_145_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_145_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_145_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_145_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_145_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_145_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_145_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_145_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_145_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_145_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_145_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_145_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_145_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_145_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_145_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_145_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_145_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_145_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_145_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_145_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_145_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_145_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_145_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_145_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_146_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_146_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_146_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_146_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_146_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_146_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_146_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_146_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_146_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_146_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_146_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_146_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_146_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_146_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_146_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_146_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_146_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_147_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_147_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_147_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_147_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_147_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_147_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_147_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_147_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_147_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_147_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_147_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_147_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_147_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_147_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_147_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_147_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_147_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_147_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_147_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_147_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_147_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_147_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_148_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_148_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_148_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_148_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_148_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_148_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_148_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_148_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_148_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_148_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_148_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_148_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_148_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_148_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_149_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_149_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_149_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_149_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_149_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_149_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_149_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_149_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_149_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_149_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_149_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_149_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_149_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_149_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_149_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_150_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_150_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_150_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_150_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_150_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_150_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_150_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_150_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_150_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_150_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_150_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_150_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_150_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_150_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_150_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_150_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_150_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_150_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_150_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_150_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_150_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_150_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_150_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_150_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_150_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_151_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_151_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_151_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_151_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_151_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_151_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_151_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_151_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_151_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_151_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_151_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_151_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_151_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_151_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_151_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_151_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_151_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_152_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_152_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_152_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_152_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_152_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_152_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_152_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_152_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_152_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_152_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_152_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_152_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_152_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_152_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_152_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_152_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_152_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_152_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_153_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_153_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_153_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_153_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_153_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_153_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_153_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_153_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_153_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_153_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_153_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_153_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_153_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_153_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_153_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_153_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_153_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_153_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_153_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_153_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_154_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_154_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_154_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_154_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_154_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_154_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_154_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_154_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_154_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_154_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_154_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_155_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_155_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_155_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_155_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_155_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_155_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_155_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_155_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_155_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_155_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_155_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_155_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_156_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_156_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_156_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_156_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_156_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_156_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_156_448 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_156_454 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_156_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_157_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_157_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_157_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_157_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_157_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_157_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_157_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_157_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_157_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_157_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_157_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_157_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_157_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_157_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_157_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_157_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_157_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_158_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_158_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_158_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_158_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_158_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_158_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_158_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_158_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_158_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_158_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_158_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_158_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_158_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_158_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_158_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_158_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_158_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_158_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_158_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_158_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_158_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_158_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_158_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_158_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_158_451 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_158_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_158_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_158_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_158_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_159_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_159_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_159_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_159_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_159_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_159_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_159_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_159_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_160_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_160_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_160_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_160_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_160_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_160_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_160_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_160_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_160_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_160_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_160_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_160_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_160_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_160_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_160_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_160_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_160_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_451 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_422 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_454 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_431 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_448 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_448 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_81_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_81_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_81_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_81_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_81_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_81_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_81_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_81_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_81_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_82_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_82_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_82_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_82_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_82_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_82_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_82_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_82_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_83_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_83_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_83_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_83_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_83_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_83_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_83_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_83_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_83_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_83_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_83_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_83_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_83_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_83_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_83_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_83_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_84_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_84_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_84_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_84_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_84_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_84_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_84_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_84_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_84_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_84_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_448 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_84_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_84_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_85_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_85_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_85_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_85_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_85_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_85_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_85_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_85_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_85_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_86_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_86_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_86_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_86_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_86_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_86_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_86_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_86_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_86_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_86_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_86_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_86_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_86_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_86_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_86_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_86_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_86_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_87_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_87_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_87_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_87_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_87_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_87_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_87_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_87_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_87_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_87_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_87_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_88_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_88_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_88_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_88_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_88_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_88_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_88_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_88_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_448 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_88_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_88_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_89_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_89_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_89_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_89_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_89_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_89_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_89_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_89_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_89_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_89_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_89_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_89_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_89_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_89_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_89_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_89_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_89_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_89_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_89_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_89_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_89_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_89_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_89_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_89_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_89_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_90_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_90_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_90_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_90_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_90_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_90_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_90_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_90_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_90_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_90_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_90_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_90_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_90_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_90_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_90_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_91_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_91_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_91_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_91_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_91_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_91_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_91_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_91_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_91_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_91_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_91_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_91_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_91_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_91_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_91_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_91_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_91_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_91_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_91_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_92_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_92_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_92_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_92_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_92_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_92_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_92_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_92_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_92_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_92_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_92_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_92_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_92_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_92_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_92_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_92_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_92_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_92_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_92_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_92_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_92_454 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_92_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_92_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_92_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_92_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_93_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_93_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_93_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_93_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_93_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_93_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_93_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_93_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_93_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_93_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_93_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_422 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_93_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_93_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_93_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_94_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_94_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_94_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_94_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_94_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_94_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_94_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_94_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_94_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_94_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_94_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_94_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_94_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_94_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_94_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_94_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_94_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_94_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_94_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_94_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_94_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_94_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_94_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_94_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_95_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_95_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_95_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_95_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_95_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_95_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_95_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_95_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_95_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_95_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_95_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_95_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_95_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_95_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_95_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_95_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_95_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_95_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_95_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_96_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_96_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_96_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_96_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_96_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_96_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_96_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_96_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_96_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_96_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_96_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_96_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_96_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_96_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_96_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_96_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_96_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_451 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_97_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_97_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_97_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_97_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_97_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_97_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_97_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_97_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_97_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_97_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_97_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_97_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_97_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_97_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_97_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_98_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_98_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_98_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_98_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_98_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_98_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_98_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_98_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_99_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_99_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_99_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_99_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_99_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_99_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_99_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_99_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_99_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_99_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_99_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_99_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_99_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_99_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_99_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_99_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_0/_0_  (.A(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_1/_0_  (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_2/_0_  (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_3/_0_  (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_4/_0_  (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_5/_0_  (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_6/_0_  (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_7/_0_  (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_8/_0_  (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_9/_0_  (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_0/_0_  (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_1/_0_  (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_10/_0_  (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_11/_0_  (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_2/_0_  (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_3/_0_  (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_4/_0_  (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_5/_0_  (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_6/_0_  (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_7/_0_  (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_8/_0_  (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_9/_0_  (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[374] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[374] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[375] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[375] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[384] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[384] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[385] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[385] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[386] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[386] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[387] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[387] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[388] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[388] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[389] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[389] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[390] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[390] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[391] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[391] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[392] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[392] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[393] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[393] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[376] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[376] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[394] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[394] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[395] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[395] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[396] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[396] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[397] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[397] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[398] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[398] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[399] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[399] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[400] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[400] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[401] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[401] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[402] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[402] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[403] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[403] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[377] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[377] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[404] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[404] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[405] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[405] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[378] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[378] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[379] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[379] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[380] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[380] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[381] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[381] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[382] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[382] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[383] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[383] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[54] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[55] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[64] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[65] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[66] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[67] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[68] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[69] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[70] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[71] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[72] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[73] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[56] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[74] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[75] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[76] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[77] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[78] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[79] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[80] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[81] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[82] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[83] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[57] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[84] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[85] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[58] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[59] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[60] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[61] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[62] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[63] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[22] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[23] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[32] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[33] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[34] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[35] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[36] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[37] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[38] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[39] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[40] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[41] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[24] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[42] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[43] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[44] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[45] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[46] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[47] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[50] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[51] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[25] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[26] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[27] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[28] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[29] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[30] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[31] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[0] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[1] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[2] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[3] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[4] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[5] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[6] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[7] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[8] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[9] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[10] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[11] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[12] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[13] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[14] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[15] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[16] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[17] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[17] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[18] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[19] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[20] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[21] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[342] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[343] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[352] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[352] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[353] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[353] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[354] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[355] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[356] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[356] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[357] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[357] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[358] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[359] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[360] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[360] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[361] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[361] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[344] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[344] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[362] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[363] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[364] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[364] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[365] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[365] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[366] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[367] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[368] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[368] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[369] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[369] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[370] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[371] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[345] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[345] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[372] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[372] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[373] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[373] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[346] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[347] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[348] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[348] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[349] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[349] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[350] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[351] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[320] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[321] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[324] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[325] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[328] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[328] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[329] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[329] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[312] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[330] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[331] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[332] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[332] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[333] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[333] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[334] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[335] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[336] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[336] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[337] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[337] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[338] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[339] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[313] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[340] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[340] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[341] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[341] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[316] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[317] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[288] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[289] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[292] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[293] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[296] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[297] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[280] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[300] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[301] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[304] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[305] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[281] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[308] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[309] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[284] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[285] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[256] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[257] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[260] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[261] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[264] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[265] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[248] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[268] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[269] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[272] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[273] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[249] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[276] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[277] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[252] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[253] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[214] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[215] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[224] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[225] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[226] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[227] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[228] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[229] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[230] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[231] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[232] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[233] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[216] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[234] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[235] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[236] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[237] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[238] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[239] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[240] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[241] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[242] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[243] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[217] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[244] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[245] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[218] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[219] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[220] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[221] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[222] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[223] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[182] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[183] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[192] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[193] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[194] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[195] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[196] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[197] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[198] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[199] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[200] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[201] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[184] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[202] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[203] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[204] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[205] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[206] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[207] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[208] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[209] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[210] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[211] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[185] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[212] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[213] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[186] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[187] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[188] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[189] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[190] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[191] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[150] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[151] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[160] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[161] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[162] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[163] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[164] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[165] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[166] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[167] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[168] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[169] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[152] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[170] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[171] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[172] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[173] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[174] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[175] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[176] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[177] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[178] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[179] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[153] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[180] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[181] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[154] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[155] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[156] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[157] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[158] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[159] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[118] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[119] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[128] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[129] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[130] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[131] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[132] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[133] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[134] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[135] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[136] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[137] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[120] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[138] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[139] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[140] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[141] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[142] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[143] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[144] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[145] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[146] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[147] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[121] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[148] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[149] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[122] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[123] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[124] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[125] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[126] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[127] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[86] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[87] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[96] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[97] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[98] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[99] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[100] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[101] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[102] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[103] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[88] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[106] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[107] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[110] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[111] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[112] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[113] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[114] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[115] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[89] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[116] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[117] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[90] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[91] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[92] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[93] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[94] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[95] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[95] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_00_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_01_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_02_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_03_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_04_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_05_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_06_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_07_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_08_  (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_09_  (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_10_  (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_11_  (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_12_  (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_13_  (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_14_  (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_15_  (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_16_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_17_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_18_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_19_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_20_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_21_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_22_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_23_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_24_  (.A(\Tile_X0Y1_N2BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_25_  (.A(\Tile_X0Y1_N2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net495));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_26_  (.A(\Tile_X0Y1_N2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_27_  (.A(\Tile_X0Y1_N2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_28_  (.A(\Tile_X0Y1_N2BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_29_  (.A(\Tile_X0Y1_N2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_30_  (.A(\Tile_X0Y1_N2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_31_  (.A(\Tile_X0Y1_N2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_32_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_33_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEG[1] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_34_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEG[2] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_35_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEG[3] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_36_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEG[4] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_37_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEG[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_38_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEG[6] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_39_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEG[7] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_40_  (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEGb[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_41_  (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEGb[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_42_  (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEGb[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_43_  (.A(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEGb[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_44_  (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEGb[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_45_  (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEGb[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_46_  (.A(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEGb[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_47_  (.A(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S2BEGb[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_48_  (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_49_  (.A(\Tile_X0Y0_DSP_top/JW2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_50_  (.A(\Tile_X0Y0_DSP_top/JW2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_51_  (.A(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_52_  (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_53_  (.A(\Tile_X0Y0_DSP_top/JW2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_54_  (.A(\Tile_X0Y0_DSP_top/JW2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_55_  (.A(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_56_  (.A(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_57_  (.A(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_58_  (.A(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_59_  (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_60_  (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_61_  (.A(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_62_  (.A(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_63_  (.A(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0  (.A0(net4),
    .A1(net136),
    .A2(\Tile_X0Y1_bot2top[0] ),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y1_bot2top[3] ),
    .A2(\Tile_X0Y1_bot2top[4] ),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y1_bot2top[7] ),
    .A2(\Tile_X0Y1_bot2top[8] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[50] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0  (.A0(net3),
    .A1(net135),
    .A2(\Tile_X0Y1_bot2top[0] ),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y1_bot2top[3] ),
    .A2(\Tile_X0Y1_bot2top[4] ),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y1_bot2top[7] ),
    .A2(\Tile_X0Y1_bot2top[8] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[54] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[1] ),
    .A2(\Tile_X0Y1_N4BEG[1] ),
    .A3(net40),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net86),
    .A2(net138),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[1] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[280] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[2] ),
    .A2(\Tile_X0Y1_N4BEG[2] ),
    .A3(net7),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net87),
    .A2(net139),
    .A3(net174),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[284] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[3] ),
    .A2(\Tile_X0Y1_N4BEG[3] ),
    .A3(net8),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net88),
    .A2(net140),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[288] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[4] ),
    .A2(\Tile_X0Y1_N4BEG[0] ),
    .A3(net9),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net89),
    .A2(net141),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[292] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[5] ),
    .A2(net2),
    .A3(net10),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net84),
    .A2(net90),
    .A3(net134),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[296] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[6] ),
    .A2(net3),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net83),
    .A2(net91),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[300] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[7] ),
    .A2(net4),
    .A3(net12),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net84),
    .A2(net92),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[304] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[0] ),
    .A2(net1),
    .A3(net5),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net83),
    .A2(net117),
    .A3(net165),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[6] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[308] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[1] ),
    .A1(\Tile_X0Y1_N4BEG[1] ),
    .A2(net4),
    .A3(net6),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net124),
    .A2(net138),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[1] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[248] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[2] ),
    .A1(\Tile_X0Y1_N4BEG[2] ),
    .A2(net1),
    .A3(net7),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net87),
    .A2(net139),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[252] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[3] ),
    .A1(\Tile_X0Y1_N4BEG[3] ),
    .A2(net2),
    .A3(net8),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net88),
    .A2(net140),
    .A3(net172),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[256] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[4] ),
    .A1(\Tile_X0Y1_N4BEG[0] ),
    .A2(net3),
    .A3(net9),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net89),
    .A2(net141),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[260] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[5] ),
    .A2(net2),
    .A3(net10),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net90),
    .A2(net134),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[264] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[6] ),
    .A2(net3),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1  (.A0(net83),
    .A1(net91),
    .A2(net133),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[268] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[7] ),
    .A2(net4),
    .A3(net12),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1  (.A0(net84),
    .A1(net92),
    .A2(net134),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[272] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[0] ),
    .A2(net1),
    .A3(net33),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net85),
    .A2(net133),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[6] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[276] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_NN4BEG[1] ),
    .A1(net4),
    .A2(net6),
    .A3(net24),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1  (.A0(net86),
    .A1(net108),
    .A2(net138),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[1] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[312] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_NN4BEG[2] ),
    .A1(net1),
    .A2(net41),
    .A3(net21),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1  (.A0(net109),
    .A1(net125),
    .A2(net139),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[316] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_NN4BEG[3] ),
    .A1(net2),
    .A2(net8),
    .A3(net24),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1  (.A0(net88),
    .A1(net110),
    .A2(net140),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[320] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[4] ),
    .A1(net3),
    .A2(net9),
    .A3(net21),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1  (.A0(net89),
    .A1(net101),
    .A2(net141),
    .A3(net173),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[324] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[5] ),
    .A2(net2),
    .A3(net10),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net90),
    .A2(net134),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[328] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[6] ),
    .A2(net3),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1  (.A0(net83),
    .A1(net91),
    .A2(net133),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[332] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[7] ),
    .A2(net4),
    .A3(net12),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1  (.A0(net84),
    .A1(net92),
    .A2(net134),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[336] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[0] ),
    .A2(net1),
    .A3(net5),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net85),
    .A2(net133),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[6] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[340] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[1] ),
    .A2(net6),
    .A3(net24),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1  (.A0(net86),
    .A1(net108),
    .A2(net138),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[1] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[344] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[2] ),
    .A2(net7),
    .A3(net21),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1  (.A0(net87),
    .A1(net109),
    .A2(net139),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[348] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[3] ),
    .A2(net8),
    .A3(net24),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1  (.A0(net88),
    .A1(net110),
    .A2(net140),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[352] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[4] ),
    .A2(net9),
    .A3(net21),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1  (.A0(net89),
    .A1(net101),
    .A2(net141),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[356] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[5] ),
    .A2(net2),
    .A3(net10),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net84),
    .A2(net90),
    .A3(net134),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[360] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[6] ),
    .A2(net3),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net83),
    .A2(net91),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[364] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[7] ),
    .A2(net4),
    .A3(net12),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net84),
    .A2(net92),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[368] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[0] ),
    .A2(net1),
    .A3(net5),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net83),
    .A2(net85),
    .A3(net133),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[6] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[372] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0  (.A0(net4),
    .A1(net136),
    .A2(\Tile_X0Y1_bot2top[0] ),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y1_bot2top[3] ),
    .A2(\Tile_X0Y1_bot2top[4] ),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y1_bot2top[7] ),
    .A2(\Tile_X0Y1_bot2top[8] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[106] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0  (.A0(net3),
    .A1(net135),
    .A2(\Tile_X0Y1_bot2top[0] ),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y1_bot2top[3] ),
    .A2(\Tile_X0Y1_bot2top[4] ),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y1_bot2top[7] ),
    .A2(\Tile_X0Y1_bot2top[8] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[110] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_E1BEG0  (.A0(\Tile_X0Y1_bot2top[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/JN2BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[28] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net382));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_E1BEG1  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/JN2BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[30] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_E1BEG2  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/JN2BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[32] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_E1BEG3  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/JN2BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[34] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0  (.A0(\Tile_X0Y1_N2BEGb[6] ),
    .A1(net11),
    .A2(net126),
    .A3(net143),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[214] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1  (.A0(\Tile_X0Y1_NN4BEG[0] ),
    .A1(net7),
    .A2(net87),
    .A3(net139),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[216] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2  (.A0(\Tile_X0Y1_N2BEGb[4] ),
    .A1(net33),
    .A2(net89),
    .A3(net141),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[218] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3  (.A0(\Tile_X0Y1_N2BEGb[0] ),
    .A1(net5),
    .A2(net85),
    .A3(net174),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[220] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0  (.A0(\Tile_X0Y1_NN4BEG[3] ),
    .A1(net11),
    .A2(net91),
    .A3(net143),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[222] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1  (.A0(\Tile_X0Y1_N2BEGb[2] ),
    .A1(net7),
    .A2(net87),
    .A3(net173),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[224] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2  (.A0(\Tile_X0Y1_N2BEGb[4] ),
    .A1(net9),
    .A2(net125),
    .A3(net141),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[226] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3  (.A0(\Tile_X0Y1_N2BEGb[0] ),
    .A1(net40),
    .A2(net85),
    .A3(net137),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[228] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0  (.A0(\Tile_X0Y1_N2BEGb[7] ),
    .A1(net41),
    .A2(net92),
    .A3(net144),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[230] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1  (.A0(\Tile_X0Y1_N2BEGb[3] ),
    .A1(net8),
    .A2(net88),
    .A3(net172),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[232] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2  (.A0(\Tile_X0Y1_N2BEGb[5] ),
    .A1(net10),
    .A2(net124),
    .A3(net142),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[234] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3  (.A0(\Tile_X0Y1_NN4BEG[2] ),
    .A1(net6),
    .A2(net86),
    .A3(net138),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[236] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0  (.A0(\Tile_X0Y1_N2BEGb[7] ),
    .A1(net12),
    .A2(net92),
    .A3(net165),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[238] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1  (.A0(\Tile_X0Y1_N2BEGb[3] ),
    .A1(net8),
    .A2(net117),
    .A3(net140),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[240] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2  (.A0(\Tile_X0Y1_NN4BEG[1] ),
    .A1(net10),
    .A2(net90),
    .A3(net142),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[242] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3  (.A0(\Tile_X0Y1_N2BEGb[1] ),
    .A1(net42),
    .A2(net86),
    .A3(net138),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[244] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2END_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0  (.A0(\Tile_X0Y1_N2BEG[6] ),
    .A1(net99),
    .A2(net151),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[150] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1  (.A0(net15),
    .A1(net95),
    .A2(net147),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[152] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2  (.A0(\Tile_X0Y1_N2BEG[4] ),
    .A1(net17),
    .A2(net149),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[154] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3  (.A0(\Tile_X0Y1_N2BEG[0] ),
    .A1(net13),
    .A2(net93),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[156] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0  (.A0(\Tile_X0Y1_N2BEG[7] ),
    .A1(net20),
    .A2(net100),
    .A3(net152),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[182] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1  (.A0(\Tile_X0Y1_N2BEG[3] ),
    .A1(net16),
    .A2(net96),
    .A3(net148),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[184] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2  (.A0(\Tile_X0Y1_N2BEG[5] ),
    .A1(net18),
    .A2(net98),
    .A3(net150),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[186] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3  (.A0(\Tile_X0Y1_N2BEG[1] ),
    .A1(net14),
    .A2(net94),
    .A3(net146),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[188] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0  (.A0(net19),
    .A1(net99),
    .A2(net151),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[158] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1  (.A0(\Tile_X0Y1_N2BEG[2] ),
    .A1(net15),
    .A2(net147),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[160] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2  (.A0(\Tile_X0Y1_N2BEG[4] ),
    .A1(net17),
    .A2(net97),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[162] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3  (.A0(\Tile_X0Y1_N2BEG[0] ),
    .A1(net93),
    .A2(net145),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[164] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0  (.A0(\Tile_X0Y1_N2BEG[7] ),
    .A1(net20),
    .A2(net100),
    .A3(net152),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[190] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1  (.A0(\Tile_X0Y1_N2BEG[3] ),
    .A1(net16),
    .A2(net96),
    .A3(net148),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[192] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2  (.A0(\Tile_X0Y1_N2BEG[5] ),
    .A1(net18),
    .A2(net98),
    .A3(net150),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[194] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3  (.A0(\Tile_X0Y1_N2BEG[1] ),
    .A1(net14),
    .A2(net94),
    .A3(net146),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[196] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0  (.A0(\Tile_X0Y1_N2BEG[6] ),
    .A1(net19),
    .A2(net151),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[166] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1  (.A0(\Tile_X0Y1_N2BEG[2] ),
    .A1(net15),
    .A2(net95),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[168] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2  (.A0(\Tile_X0Y1_N2BEG[4] ),
    .A1(net97),
    .A2(net149),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[170] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3  (.A0(net13),
    .A1(net93),
    .A2(net145),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[172] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0  (.A0(\Tile_X0Y1_N2BEG[7] ),
    .A1(net20),
    .A2(net100),
    .A3(net152),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[198] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1  (.A0(\Tile_X0Y1_N2BEG[3] ),
    .A1(net16),
    .A2(net96),
    .A3(net148),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[200] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2  (.A0(\Tile_X0Y1_N2BEG[5] ),
    .A1(net18),
    .A2(net98),
    .A3(net150),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[202] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3  (.A0(\Tile_X0Y1_N2BEG[1] ),
    .A1(net14),
    .A2(net94),
    .A3(net146),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[204] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0  (.A0(\Tile_X0Y1_N2BEG[6] ),
    .A1(net19),
    .A2(net99),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[174] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1  (.A0(\Tile_X0Y1_N2BEG[2] ),
    .A1(net95),
    .A2(net147),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[176] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2  (.A0(net17),
    .A1(net97),
    .A2(net149),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[178] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3  (.A0(\Tile_X0Y1_N2BEG[0] ),
    .A1(net13),
    .A2(net145),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[180] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0  (.A0(\Tile_X0Y1_N2BEG[7] ),
    .A1(net20),
    .A2(net100),
    .A3(net152),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[206] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1  (.A0(\Tile_X0Y1_N2BEG[3] ),
    .A1(net16),
    .A2(net96),
    .A3(net148),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[208] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2  (.A0(\Tile_X0Y1_N2BEG[5] ),
    .A1(net18),
    .A2(net98),
    .A3(net150),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[210] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3  (.A0(\Tile_X0Y1_N2BEG[1] ),
    .A1(net14),
    .A2(net94),
    .A3(net146),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[212] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0  (.A0(\Tile_X0Y1_NN4BEG[3] ),
    .A1(net110),
    .A2(net165),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[374] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[375] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1  (.A0(net41),
    .A1(net109),
    .A2(net144),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[376] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2  (.A0(\Tile_X0Y1_N4BEG[1] ),
    .A1(net24),
    .A2(net156),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[378] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[379] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3  (.A0(\Tile_X0Y1_N4BEG[0] ),
    .A1(net21),
    .A2(net101),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[380] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0  (.A0(net8),
    .A1(net126),
    .A2(net173),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[382] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[383] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1  (.A0(\Tile_X0Y1_N4BEG[2] ),
    .A1(net7),
    .A2(net144),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[384] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[385] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2  (.A0(\Tile_X0Y1_NN4BEG[1] ),
    .A1(net40),
    .A2(net108),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[386] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[387] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3  (.A0(\Tile_X0Y1_N4BEG[0] ),
    .A1(net117),
    .A2(net153),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[388] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[389] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0  (.A0(\Tile_X0Y1_N4BEG[3] ),
    .A1(net8),
    .A2(net140),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[390] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[391] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1  (.A0(\Tile_X0Y1_NN4BEG[2] ),
    .A1(net7),
    .A2(net109),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[392] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[393] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2  (.A0(\Tile_X0Y1_N4BEG[1] ),
    .A1(net124),
    .A2(net141),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[394] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[395] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3  (.A0(net42),
    .A1(net101),
    .A2(net172),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[396] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[397] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0  (.A0(\Tile_X0Y1_N4BEG[3] ),
    .A1(net33),
    .A2(net110),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[398] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[399] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1  (.A0(\Tile_X0Y1_N4BEG[2] ),
    .A1(net125),
    .A2(net139),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[400] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[401] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2  (.A0(net24),
    .A1(net108),
    .A2(net174),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[402] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[403] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3  (.A0(\Tile_X0Y1_NN4BEG[0] ),
    .A1(net21),
    .A2(net137),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[404] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[405] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N1BEG0  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[0] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N1BEG1  (.A0(\Tile_X0Y1_bot2top[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[2] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net483));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N1BEG2  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[4] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net484));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N1BEG3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[6] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net485));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N4BEG0  (.A0(\Tile_X0Y1_N2BEGb[2] ),
    .A1(\Tile_X0Y1_N4BEG[1] ),
    .A2(net24),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[8] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N4BEG1  (.A0(\Tile_X0Y1_N2BEGb[3] ),
    .A1(\Tile_X0Y1_N4BEG[2] ),
    .A2(net21),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[10] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N4BEG2  (.A0(\Tile_X0Y1_N2BEGb[0] ),
    .A1(\Tile_X0Y1_N4BEG[3] ),
    .A2(net156),
    .A3(\Tile_X0Y1_bot2top[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[12] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net507));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N4BEG3  (.A0(\Tile_X0Y1_N2BEGb[1] ),
    .A1(\Tile_X0Y1_N4BEG[0] ),
    .A2(net153),
    .A3(\Tile_X0Y1_bot2top[7] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[14] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net508));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S1BEG0  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[56] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S1BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S1BEG1  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[58] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S1BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S1BEG2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[60] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S1BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S1BEG3  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[62] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S1BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S4BEG0  (.A0(net24),
    .A1(net87),
    .A2(net108),
    .A3(\Tile_X0Y1_bot2top[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[64] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S4BEG1  (.A0(net21),
    .A1(net88),
    .A2(net109),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[66] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S4BEG2  (.A0(net85),
    .A1(net110),
    .A2(net156),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[68] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S4BEG3  (.A0(net86),
    .A1(net101),
    .A2(net153),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[70] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_W1BEG0  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/JS2BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[84] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_W1BEG1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/JS2BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[86] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_W1BEG2  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/JS2BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[88] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_W1BEG3  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/JS2BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[90] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot0  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_AB_BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[112] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot1  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_AB_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[114] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot10  (.A0(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_EF_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[132] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[10] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot11  (.A0(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_EF_BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[134] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[11] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot12  (.A0(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_GH_BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[136] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot13  (.A0(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_GH_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[138] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot14  (.A0(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[140] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot15  (.A0(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_GH_BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[142] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot2  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_AB_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[116] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_AB_BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[118] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot4  (.A0(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_CD_BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[120] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot5  (.A0(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_CD_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[122] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot6  (.A0(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_CD_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[124] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot7  (.A0(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_CD_BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[126] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[7] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot8  (.A0(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_EF_BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[128] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[8] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot9  (.A0(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_EF_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[130] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_top2bot[9] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(net3),
    .A2(net83),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[36] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_GH_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[36] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[38] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net417));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(net4),
    .A2(net84),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[39] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_EF_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[39] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[41] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net418));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(net1),
    .A2(net81),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[42] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[8] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_CD_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[42] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[44] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net419));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(net2),
    .A2(net82),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[45] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[9] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[45] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[47] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net420));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(net3),
    .A2(net135),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[16] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_GH_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[16] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[18] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net521));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(net4),
    .A2(net136),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[19] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_EF_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[19] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[21] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net522));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(net1),
    .A2(net133),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[22] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[8] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[22] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[24] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net523));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(net2),
    .A2(net134),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[25] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[9] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_AB_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[25] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[27] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net524));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(net3),
    .A2(net135),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[72] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[72] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[74] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_SS4BEG[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(net4),
    .A2(net136),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[75] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_EF_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[75] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[77] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_SS4BEG[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(net1),
    .A2(net133),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[78] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[8] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_CD_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[78] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[80] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_SS4BEG[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(net2),
    .A2(net134),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[81] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[9] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_AB_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[81] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[83] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_SS4BEG[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(net83),
    .A2(net135),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[92] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[92] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[94] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net570));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(net84),
    .A2(net136),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[95] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[95] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[97] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net571));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(net81),
    .A2(net133),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[98] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[8] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_CD_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[98] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[100] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net572));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(net82),
    .A2(net134),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[101] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[9] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_AB_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[101] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[103] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net573));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_inst0  (.A0(\Tile_X0Y0_DSP_top/JN2BEG[4] ),
    .A1(\Tile_X0Y0_DSP_top/JN2BEG[6] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[4] ),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[144] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_DSP_top/JS2BEG[4] ),
    .A1(\Tile_X0Y0_DSP_top/JS2BEG[6] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[4] ),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[144] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[146] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_top2bot[16] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_inst0  (.A0(\Tile_X0Y0_DSP_top/JN2BEG[5] ),
    .A1(\Tile_X0Y0_DSP_top/JN2BEG[7] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[5] ),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[7] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[147] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_DSP_top/JS2BEG[5] ),
    .A1(\Tile_X0Y0_DSP_top/JS2BEG[7] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[5] ),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[7] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[147] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[149] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y0_top2bot[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net517));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_0/_0_  (.A(\Tile_X0Y1_N4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[0] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_1/_0_  (.A(\Tile_X0Y1_N4BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/N4END_inbuf_10/_0_  (.A(\Tile_X0Y1_N4BEG[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/N4END_inbuf_11/_0_  (.A(\Tile_X0Y1_N4BEG[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[11] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_2/_0_  (.A(\Tile_X0Y1_N4BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_3/_0_  (.A(\Tile_X0Y1_N4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[3] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_4/_0_  (.A(\Tile_X0Y1_N4BEG[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_5/_0_  (.A(\Tile_X0Y1_N4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[5] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_6/_0_  (.A(\Tile_X0Y1_N4BEG[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[6] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_7/_0_  (.A(\Tile_X0Y1_N4BEG[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/N4END_inbuf_8/_0_  (.A(\Tile_X0Y1_N4BEG[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[8] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_9/_0_  (.A(\Tile_X0Y1_N4BEG[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_0/_0_  (.A(\Tile_X0Y1_NN4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[0] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_1/_0_  (.A(\Tile_X0Y1_NN4BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_10/_0_  (.A(\Tile_X0Y1_NN4BEG[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_11/_0_  (.A(\Tile_X0Y1_NN4BEG[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_2/_0_  (.A(\Tile_X0Y1_NN4BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_3/_0_  (.A(\Tile_X0Y1_NN4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_4/_0_  (.A(\Tile_X0Y1_NN4BEG[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_5/_0_  (.A(\Tile_X0Y1_NN4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_6/_0_  (.A(\Tile_X0Y1_NN4BEG[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_7/_0_  (.A(\Tile_X0Y1_NN4BEG[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_8/_0_  (.A(\Tile_X0Y1_NN4BEG[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[8] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_9/_0_  (.A(\Tile_X0Y1_NN4BEG[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[9] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/S4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_S4BEG[9] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_0/_0_  (.A(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_1/_0_  (.A(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_10/_0_  (.A(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_11/_0_  (.A(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_2/_0_  (.A(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[2] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_3/_0_  (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_4/_0_  (.A(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[4] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/S4END_inbuf_5/_0_  (.A(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_6/_0_  (.A(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_7/_0_  (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_8/_0_  (.A(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_9/_0_  (.A(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[10] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[11] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[3] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[4] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[6] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[8] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_SS4BEG[9] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4END_inbuf_0/_0_  (.A(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/SS4END_inbuf_1/_0_  (.A(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_10/_0_  (.A(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_11/_0_  (.A(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4END_inbuf_2/_0_  (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[2] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/SS4END_inbuf_3/_0_  (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_4/_0_  (.A(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_5/_0_  (.A(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_6/_0_  (.A(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_7/_0_  (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_8/_0_  (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_9/_0_  (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_0/_0_  (.A(net157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_1/_0_  (.A(net158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_2/_0_  (.A(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_3/_0_  (.A(net160),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_4/_0_  (.A(net161),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_5/_0_  (.A(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_6/_0_  (.A(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_7/_0_  (.A(net164),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_8/_0_  (.A(net154),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_9/_0_  (.A(net155),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_0/_0_  (.A(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_1/_0_  (.A(net176),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_10/_0_  (.A(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_11/_0_  (.A(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_2/_0_  (.A(net177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_3/_0_  (.A(net178),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_4/_0_  (.A(net179),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_5/_0_  (.A(net180),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_6/_0_  (.A(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_7/_0_  (.A(net167),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_8/_0_  (.A(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_9/_0_  (.A(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_0/_0_  (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_1/_0_  (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_10/_0_  (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_11/_0_  (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_12/_0_  (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_13/_0_  (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_14/_0_  (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_15/_0_  (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_16/_0_  (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[16] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/data_inbuf_17/_0_  (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_18/_0_  (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_19/_0_  (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_2/_0_  (.A(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_20/_0_  (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[20] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_21/_0_  (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[21] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_22/_0_  (.A(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[22] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_23/_0_  (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[23] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_24/_0_  (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[24] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_25/_0_  (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[25] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_26/_0_  (.A(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[26] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_27/_0_  (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[27] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_28/_0_  (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[28] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_29/_0_  (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[29] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_3/_0_  (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[3] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/data_inbuf_30/_0_  (.A(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[30] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/data_inbuf_31/_0_  (.A(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[31] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_4/_0_  (.A(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_5/_0_  (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_6/_0_  (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_7/_0_  (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_8/_0_  (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_9/_0_  (.A(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_12/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_13/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_14/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_15/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_16/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_17/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_18/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_19/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_20/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_21/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_22/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_23/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_24/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_25/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_26/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_27/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_28/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_29/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_30/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_31/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/inst_clk_buf  (.A(Tile_X0Y1_UserCLKo),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_0/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_1/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_10/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_11/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_12/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_13/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_14/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_15/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_16/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_17/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_18/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_19/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_2/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_3/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_4/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_5/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_6/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_7/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_8/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_9/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[9] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net462));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net464));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_12/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_13/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_14/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_15/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_16/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_17/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_18/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_19/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net472));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net477));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net480));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_0/_0_  (.A(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_1/_0_  (.A(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_2/_0_  (.A(net207),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_3/_0_  (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_4/_0_  (.A(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_5/_0_  (.A(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_6/_0_  (.A(net211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_7/_0_  (.A(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_8/_0_  (.A(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_9/_0_  (.A(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_0/_0_  (.A(net223),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_1/_0_  (.A(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_10/_0_  (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_11/_0_  (.A(net219),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_2/_0_  (.A(net225),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_3/_0_  (.A(net226),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_4/_0_  (.A(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_5/_0_  (.A(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_6/_0_  (.A(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_7/_0_  (.A(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_8/_0_  (.A(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_9/_0_  (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit0  (.D(net229),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[384] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[384] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit1  (.D(net240),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[385] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[385] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit10  (.D(net230),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[394] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[394] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit11  (.D(net231),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[395] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[395] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit12  (.D(net232),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[396] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[396] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit13  (.D(net233),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[397] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[397] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit14  (.D(net234),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[398] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[398] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit15  (.D(net235),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[399] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[399] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit16  (.D(net236),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[400] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[400] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit17  (.D(net237),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[401] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[401] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit18  (.D(net238),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[402] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[402] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit19  (.D(net239),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[403] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[403] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit2  (.D(net251),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[386] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[386] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit20  (.D(net241),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[404] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[404] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit21  (.D(net242),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[405] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[405] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit22  (.D(net243),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[406] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[406] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit23  (.D(net244),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[407] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[407] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit24  (.D(net245),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[408] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[408] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit25  (.D(net246),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[409] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[409] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit26  (.D(net247),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[410] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[410] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit27  (.D(net248),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[411] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[411] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit28  (.D(net249),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[412] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[412] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit29  (.D(net250),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[413] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[413] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit3  (.D(net254),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[387] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[387] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit30  (.D(net252),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[414] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[414] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit31  (.D(net253),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[415] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[415] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit4  (.D(net255),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[388] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[388] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit5  (.D(net256),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[389] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[389] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit6  (.D(net257),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[390] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[390] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit7  (.D(net258),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[391] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[391] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit8  (.D(net259),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[392] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[392] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit9  (.D(net260),
    .GATE(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[393] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[393] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit0  (.D(net229),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[64] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit1  (.D(net240),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[65] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit10  (.D(net230),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[74] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit11  (.D(net231),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[75] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit12  (.D(net232),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[76] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit13  (.D(net233),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[77] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit14  (.D(net234),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[78] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit15  (.D(net235),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[79] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit16  (.D(net236),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[80] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit17  (.D(net237),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[81] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit18  (.D(net238),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[82] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit19  (.D(net239),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[83] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit2  (.D(net251),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[66] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit20  (.D(net241),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[84] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit21  (.D(net242),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[85] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit22  (.D(net243),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[86] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit23  (.D(net244),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[87] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit24  (.D(net245),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[88] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit25  (.D(net246),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[89] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit26  (.D(net247),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[90] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit27  (.D(net248),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[91] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit28  (.D(net249),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[92] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit29  (.D(net250),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[93] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit3  (.D(net254),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[67] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit30  (.D(net252),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[94] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit31  (.D(net253),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[95] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit4  (.D(net255),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[68] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit5  (.D(net256),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[69] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit6  (.D(net257),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[70] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit7  (.D(net258),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[71] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit8  (.D(net259),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[72] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit9  (.D(net260),
    .GATE(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[73] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit0  (.D(net229),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[32] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit1  (.D(net240),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[33] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit10  (.D(net230),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[42] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit11  (.D(net231),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[43] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit12  (.D(net232),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[44] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit13  (.D(net233),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[45] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit14  (.D(net234),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[46] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit15  (.D(net235),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[47] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit16  (.D(net236),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[48] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit17  (.D(net237),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[49] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit18  (.D(net238),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[50] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit19  (.D(net239),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[51] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit2  (.D(net251),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[34] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit20  (.D(net241),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[52] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit21  (.D(net242),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[53] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit22  (.D(net243),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit23  (.D(net244),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit24  (.D(net245),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[56] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit25  (.D(net246),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[57] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit26  (.D(net247),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit27  (.D(net248),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit28  (.D(net249),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[60] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit29  (.D(net250),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[61] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit3  (.D(net254),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[35] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit30  (.D(net252),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[62] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit31  (.D(net253),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[63] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit4  (.D(net255),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[36] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit5  (.D(net256),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[37] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit6  (.D(net257),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[38] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit7  (.D(net258),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[39] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit8  (.D(net259),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[40] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit9  (.D(net260),
    .GATE(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[41] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit0  (.D(net229),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[0] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit1  (.D(net240),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit10  (.D(net230),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[10] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit11  (.D(net231),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[11] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit12  (.D(net232),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[12] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit13  (.D(net233),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[13] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit14  (.D(net234),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[14] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit15  (.D(net235),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[15] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit16  (.D(net236),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[16] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit17  (.D(net237),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[17] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[17] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit18  (.D(net238),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[18] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit19  (.D(net239),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[19] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit2  (.D(net251),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[2] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit20  (.D(net241),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[20] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit21  (.D(net242),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[21] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit22  (.D(net243),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[22] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit23  (.D(net244),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[23] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit24  (.D(net245),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[24] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit25  (.D(net246),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[25] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit26  (.D(net247),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[26] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit27  (.D(net248),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[27] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit28  (.D(net249),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[28] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit29  (.D(net250),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[29] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit3  (.D(net254),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[3] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit30  (.D(net252),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[30] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit31  (.D(net253),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[31] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit4  (.D(net255),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit5  (.D(net256),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit6  (.D(net257),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[6] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit7  (.D(net258),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[7] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit8  (.D(net259),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[8] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit9  (.D(net260),
    .GATE(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[9] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit0  (.D(net229),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[352] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit1  (.D(net240),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[353] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit10  (.D(net230),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[362] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[362] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit11  (.D(net231),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[363] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[363] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit12  (.D(net232),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[364] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit13  (.D(net233),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[365] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit14  (.D(net234),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[366] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[366] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit15  (.D(net235),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[367] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[367] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit16  (.D(net236),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[368] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit17  (.D(net237),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[369] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit18  (.D(net238),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[370] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[370] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit19  (.D(net239),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[371] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[371] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit2  (.D(net251),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[354] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[354] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit20  (.D(net241),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[372] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit21  (.D(net242),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[373] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit22  (.D(net243),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[374] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[374] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit23  (.D(net244),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[375] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[375] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit24  (.D(net245),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[376] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit25  (.D(net246),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[377] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit26  (.D(net247),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[378] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[378] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit27  (.D(net248),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[379] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[379] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit28  (.D(net249),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[380] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit29  (.D(net250),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[381] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit3  (.D(net254),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[355] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[355] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit30  (.D(net252),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[382] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[382] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit31  (.D(net253),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[383] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[383] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit4  (.D(net255),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[356] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit5  (.D(net256),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[357] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit6  (.D(net257),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[358] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[358] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit7  (.D(net258),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[359] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[359] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit8  (.D(net259),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[360] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit9  (.D(net260),
    .GATE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[361] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit0  (.D(net229),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit1  (.D(net240),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit10  (.D(net230),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[330] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[330] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit11  (.D(net231),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[331] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[331] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit12  (.D(net232),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[332] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit13  (.D(net233),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[333] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit14  (.D(net234),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[334] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[334] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit15  (.D(net235),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[335] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[335] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit16  (.D(net236),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[336] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit17  (.D(net237),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[337] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit18  (.D(net238),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[338] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[338] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit19  (.D(net239),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[339] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[339] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit2  (.D(net251),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[322] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit20  (.D(net241),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[340] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit21  (.D(net242),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[341] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit22  (.D(net243),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[342] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[342] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit23  (.D(net244),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[343] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[343] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit24  (.D(net245),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[344] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit25  (.D(net246),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[345] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit26  (.D(net247),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[346] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[346] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit27  (.D(net248),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[347] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[347] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit28  (.D(net249),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[348] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit29  (.D(net250),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[349] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit3  (.D(net254),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[323] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit30  (.D(net252),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[350] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[350] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit31  (.D(net253),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[351] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[351] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit4  (.D(net255),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit5  (.D(net256),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit6  (.D(net257),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[326] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit7  (.D(net258),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[327] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit8  (.D(net259),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[328] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit9  (.D(net260),
    .GATE(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[329] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit0  (.D(net229),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit1  (.D(net240),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit10  (.D(net230),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[298] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit11  (.D(net231),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[299] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit12  (.D(net232),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit13  (.D(net233),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit14  (.D(net234),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[302] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit15  (.D(net235),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[303] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit16  (.D(net236),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit17  (.D(net237),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit18  (.D(net238),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[306] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit19  (.D(net239),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[307] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit2  (.D(net251),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[290] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit20  (.D(net241),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit21  (.D(net242),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit22  (.D(net243),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[310] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit23  (.D(net244),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[311] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit24  (.D(net245),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit25  (.D(net246),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit26  (.D(net247),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[314] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit27  (.D(net248),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[315] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit28  (.D(net249),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit29  (.D(net250),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit3  (.D(net254),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[291] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit30  (.D(net252),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[318] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit31  (.D(net253),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[319] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit4  (.D(net255),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit5  (.D(net256),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit6  (.D(net257),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[294] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit7  (.D(net258),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[295] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit8  (.D(net259),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit9  (.D(net260),
    .GATE(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit0  (.D(net229),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit1  (.D(net240),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit10  (.D(net230),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[266] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit11  (.D(net231),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[267] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit12  (.D(net232),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit13  (.D(net233),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit14  (.D(net234),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[270] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit15  (.D(net235),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[271] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit16  (.D(net236),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit17  (.D(net237),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit18  (.D(net238),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[274] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit19  (.D(net239),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[275] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit2  (.D(net251),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[258] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit20  (.D(net241),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit21  (.D(net242),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit22  (.D(net243),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[278] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit23  (.D(net244),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[279] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit24  (.D(net245),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit25  (.D(net246),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit26  (.D(net247),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[282] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit27  (.D(net248),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[283] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit28  (.D(net249),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit29  (.D(net250),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit3  (.D(net254),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[259] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit30  (.D(net252),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[286] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit31  (.D(net253),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[287] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit4  (.D(net255),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit5  (.D(net256),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit6  (.D(net257),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[262] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit7  (.D(net258),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[263] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit8  (.D(net259),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit9  (.D(net260),
    .GATE(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit0  (.D(net229),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[224] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit1  (.D(net240),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[225] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit10  (.D(net230),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[234] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit11  (.D(net231),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[235] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit12  (.D(net232),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[236] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit13  (.D(net233),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[237] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit14  (.D(net234),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[238] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit15  (.D(net235),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[239] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit16  (.D(net236),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[240] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit17  (.D(net237),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[241] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit18  (.D(net238),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[242] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit19  (.D(net239),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[243] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit2  (.D(net251),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[226] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit20  (.D(net241),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[244] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit21  (.D(net242),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[245] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit22  (.D(net243),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[246] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit23  (.D(net244),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[247] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit24  (.D(net245),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[248] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit25  (.D(net246),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[249] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit26  (.D(net247),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[250] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit27  (.D(net248),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[251] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit28  (.D(net249),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[252] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit29  (.D(net250),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[253] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit3  (.D(net254),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[227] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit30  (.D(net252),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[254] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit31  (.D(net253),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[255] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit4  (.D(net255),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[228] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit5  (.D(net256),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[229] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit6  (.D(net257),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[230] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit7  (.D(net258),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[231] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit8  (.D(net259),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[232] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit9  (.D(net260),
    .GATE(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[233] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit0  (.D(net229),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[192] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit1  (.D(net240),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[193] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit10  (.D(net230),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[202] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit11  (.D(net231),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[203] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit12  (.D(net232),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[204] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit13  (.D(net233),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[205] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit14  (.D(net234),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[206] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit15  (.D(net235),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[207] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit16  (.D(net236),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[208] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit17  (.D(net237),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[209] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit18  (.D(net238),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[210] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit19  (.D(net239),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[211] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit2  (.D(net251),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[194] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit20  (.D(net241),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[212] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit21  (.D(net242),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[213] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit22  (.D(net243),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[214] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit23  (.D(net244),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[215] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit24  (.D(net245),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[216] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit25  (.D(net246),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[217] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit26  (.D(net247),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[218] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit27  (.D(net248),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[219] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit28  (.D(net249),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[220] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit29  (.D(net250),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[221] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit3  (.D(net254),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[195] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit30  (.D(net252),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[222] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit31  (.D(net253),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[223] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit4  (.D(net255),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[196] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit5  (.D(net256),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[197] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit6  (.D(net257),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[198] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit7  (.D(net258),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[199] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit8  (.D(net259),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[200] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit9  (.D(net260),
    .GATE(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[201] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit0  (.D(net229),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[160] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit1  (.D(net240),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[161] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit10  (.D(net230),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[170] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit11  (.D(net231),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[171] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit12  (.D(net232),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[172] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit13  (.D(net233),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[173] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit14  (.D(net234),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[174] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit15  (.D(net235),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[175] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit16  (.D(net236),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[176] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit17  (.D(net237),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[177] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit18  (.D(net238),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[178] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit19  (.D(net239),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[179] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit2  (.D(net251),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[162] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit20  (.D(net241),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[180] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit21  (.D(net242),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[181] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit22  (.D(net243),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[182] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit23  (.D(net244),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[183] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit24  (.D(net245),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[184] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit25  (.D(net246),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[185] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit26  (.D(net247),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[186] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit27  (.D(net248),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[187] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit28  (.D(net249),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[188] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit29  (.D(net250),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[189] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit3  (.D(net254),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[163] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit30  (.D(net252),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[190] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit31  (.D(net253),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[191] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit4  (.D(net255),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[164] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit5  (.D(net256),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[165] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit6  (.D(net257),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[166] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit7  (.D(net258),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[167] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit8  (.D(net259),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[168] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit9  (.D(net260),
    .GATE(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[169] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit0  (.D(net229),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[128] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit1  (.D(net240),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[129] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit10  (.D(net230),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[138] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit11  (.D(net231),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[139] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit12  (.D(net232),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[140] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit13  (.D(net233),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[141] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit14  (.D(net234),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[142] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit15  (.D(net235),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[143] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit16  (.D(net236),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[144] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit17  (.D(net237),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[145] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit18  (.D(net238),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[146] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit19  (.D(net239),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[147] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit2  (.D(net251),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[130] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit20  (.D(net241),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[148] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit21  (.D(net242),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[149] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit22  (.D(net243),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[150] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit23  (.D(net244),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[151] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit24  (.D(net245),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[152] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit25  (.D(net246),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[153] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit26  (.D(net247),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[154] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit27  (.D(net248),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[155] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit28  (.D(net249),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit29  (.D(net250),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit3  (.D(net254),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[131] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit30  (.D(net252),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[158] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit31  (.D(net253),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[159] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit4  (.D(net255),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[132] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit5  (.D(net256),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[133] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit6  (.D(net257),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[134] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit7  (.D(net258),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[135] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit8  (.D(net259),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[136] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit9  (.D(net260),
    .GATE(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[137] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit0  (.D(net229),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[96] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit1  (.D(net240),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[97] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit10  (.D(net230),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[106] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit11  (.D(net231),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[107] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit12  (.D(net232),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[108] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit13  (.D(net233),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[109] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit14  (.D(net234),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit15  (.D(net235),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit16  (.D(net236),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[112] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit17  (.D(net237),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[113] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit18  (.D(net238),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit19  (.D(net239),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit2  (.D(net251),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[98] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit20  (.D(net241),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[116] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit21  (.D(net242),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[117] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit22  (.D(net243),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[118] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit23  (.D(net244),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[119] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit24  (.D(net245),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[120] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit25  (.D(net246),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[121] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit26  (.D(net247),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[122] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit27  (.D(net248),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[123] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit28  (.D(net249),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[124] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit29  (.D(net250),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[125] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit3  (.D(net254),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[99] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit30  (.D(net252),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[126] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit31  (.D(net253),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[127] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit4  (.D(net255),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[100] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit5  (.D(net256),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[101] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit6  (.D(net257),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[102] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit7  (.D(net258),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[103] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit8  (.D(net259),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[104] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit9  (.D(net260),
    .GATE(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[105] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[105] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_04_  (.A(\Tile_X0Y0_top2bot[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/A4 ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_05_  (.A(\Tile_X0Y0_top2bot[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/A5 ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_06_  (.A(\Tile_X0Y0_top2bot[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/A6 ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_07_  (.A(\Tile_X0Y0_top2bot[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/A7 ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_08_  (.A(\Tile_X0Y0_top2bot[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/B4 ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_09_  (.A(\Tile_X0Y0_top2bot[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/B5 ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_10_  (.A(\Tile_X0Y0_top2bot[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/B6 ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_11_  (.A(\Tile_X0Y0_top2bot[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/B7 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_12_  (.A(\Tile_X0Y0_top2bot[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C10 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_13_  (.A(\Tile_X0Y0_top2bot[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C11 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_14_  (.A(\Tile_X0Y0_top2bot[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C12 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_15_  (.A(\Tile_X0Y0_top2bot[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C13 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_16_  (.A(\Tile_X0Y0_top2bot[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C14 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_17_  (.A(\Tile_X0Y0_top2bot[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C15 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_18_  (.A(\Tile_X0Y0_top2bot[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C16 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_19_  (.A(\Tile_X0Y0_top2bot[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C17 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_20_  (.A(\Tile_X0Y0_top2bot[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C18 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_21_  (.A(\Tile_X0Y0_top2bot[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C19 ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_22_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_23_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_24_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_25_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_26_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_27_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_28_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_29_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_30_  (.A(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_31_  (.A(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_32_  (.A(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_33_  (.A(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_34_  (.A(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_35_  (.A(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_36_  (.A(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_37_  (.A(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_38_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_39_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEG[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_40_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEG[2] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_41_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEG[3] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_42_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEG[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_43_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEG[5] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_44_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEG[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_45_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEG[7] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_46_  (.A(net293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEGb[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_47_  (.A(net294),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEGb[1] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_48_  (.A(net295),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEGb[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_49_  (.A(net296),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEGb[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_50_  (.A(net297),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEGb[4] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_51_  (.A(net298),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEGb[5] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_52_  (.A(net299),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEGb[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_53_  (.A(net300),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N2BEGb[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_54_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_55_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_56_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_57_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_58_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_59_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_60_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_61_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_62_  (.A(\Tile_X0Y0_S2BEG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_63_  (.A(\Tile_X0Y0_S2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_64_  (.A(\Tile_X0Y0_S2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_65_  (.A(\Tile_X0Y0_S2BEG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_66_  (.A(\Tile_X0Y0_S2BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_67_  (.A(\Tile_X0Y0_S2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_68_  (.A(\Tile_X0Y0_S2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_69_  (.A(\Tile_X0Y0_S2BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_70_  (.A(net338),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_71_  (.A(\Tile_X0Y1_DSP_bot/JW2BEG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net720));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_72_  (.A(\Tile_X0Y1_DSP_bot/JW2BEG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_73_  (.A(net341),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_74_  (.A(net342),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_75_  (.A(\Tile_X0Y1_DSP_bot/JW2BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_76_  (.A(\Tile_X0Y1_DSP_bot/JW2BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_77_  (.A(net345),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_78_  (.A(net346),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net727));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_79_  (.A(net347),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_80_  (.A(net348),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_81_  (.A(net349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_82_  (.A(net350),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_83_  (.A(net351),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_84_  (.A(net352),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_85_  (.A(net353),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net734));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_86_  (.A(\Tile_X0Y1_DSP_bot/Q10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[0] ));
 sky130_fd_sc_hd__clkbuf_16 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_87_  (.A(\Tile_X0Y1_DSP_bot/Q11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[1] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_88_  (.A(\Tile_X0Y1_DSP_bot/Q12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[2] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_89_  (.A(\Tile_X0Y1_DSP_bot/Q13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[3] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_90_  (.A(\Tile_X0Y1_DSP_bot/Q14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[4] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_91_  (.A(\Tile_X0Y1_DSP_bot/Q15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[5] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_92_  (.A(\Tile_X0Y1_DSP_bot/Q16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[6] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_93_  (.A(\Tile_X0Y1_DSP_bot/Q17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[7] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_94_  (.A(\Tile_X0Y1_DSP_bot/Q18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[8] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_95_  (.A(\Tile_X0Y1_DSP_bot/Q19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_bot2top[9] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0  (.A0(net184),
    .A1(net337),
    .A2(\Tile_X0Y1_DSP_bot/Q0 ),
    .A3(\Tile_X0Y1_DSP_bot/Q1 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/Q3 ),
    .A2(\Tile_X0Y1_DSP_bot/Q4 ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/Q7 ),
    .A2(\Tile_X0Y1_DSP_bot/Q8 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[56] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0  (.A0(net183),
    .A1(net336),
    .A2(\Tile_X0Y1_DSP_bot/Q0 ),
    .A3(\Tile_X0Y1_DSP_bot/Q1 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/Q3 ),
    .A2(\Tile_X0Y1_DSP_bot/Q4 ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/Q7 ),
    .A2(\Tile_X0Y1_DSP_bot/Q8 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[60] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net286),
    .A2(net308),
    .A3(net220),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1  (.A0(net204),
    .A1(\Tile_X0Y0_S2BEGb[1] ),
    .A2(net339),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q1 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[290] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net287),
    .A2(net309),
    .A3(net187),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[2] ),
    .A2(net340),
    .A3(net375),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[294] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net288),
    .A2(net310),
    .A3(net188),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1  (.A0(net204),
    .A1(\Tile_X0Y0_S2BEGb[3] ),
    .A2(net341),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[298] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net289),
    .A2(net301),
    .A3(net189),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[4] ),
    .A2(net342),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[302] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net290),
    .A2(net182),
    .A3(net190),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(\Tile_X0Y0_S2BEGb[5] ),
    .A3(net335),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[306] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net291),
    .A2(net183),
    .A3(net191),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(\Tile_X0Y0_S2BEGb[6] ),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[310] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net292),
    .A2(net184),
    .A3(net192),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(\Tile_X0Y0_S2BEGb[7] ),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[314] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net285),
    .A2(net181),
    .A3(net185),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(\Tile_X0Y0_SS4BEG[0] ),
    .A3(net366),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(net763),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[318] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0  (.A0(net286),
    .A1(net308),
    .A2(net184),
    .A3(net186),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1  (.A0(net204),
    .A1(\Tile_X0Y0_SS4BEG[1] ),
    .A2(net339),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2  (.A0(net764),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[258] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0  (.A0(net287),
    .A1(net309),
    .A2(net181),
    .A3(net187),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[2] ),
    .A2(net340),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[262] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0  (.A0(net288),
    .A1(net310),
    .A2(net182),
    .A3(net188),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1  (.A0(net204),
    .A1(\Tile_X0Y0_S2BEGb[3] ),
    .A2(net341),
    .A3(net373),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[266] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0  (.A0(net289),
    .A1(net301),
    .A2(net183),
    .A3(net189),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[4] ),
    .A2(net342),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[270] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net290),
    .A2(net182),
    .A3(net190),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S2BEGb[5] ),
    .A2(net335),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[274] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net291),
    .A2(net183),
    .A3(net191),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[2] ),
    .A1(\Tile_X0Y0_S2BEGb[6] ),
    .A2(net334),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[278] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net292),
    .A2(net184),
    .A3(net192),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[3] ),
    .A1(\Tile_X0Y0_S2BEGb[7] ),
    .A2(net335),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[282] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net285),
    .A2(net181),
    .A3(net213),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S2BEGb[0] ),
    .A2(net334),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(net763),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[286] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0  (.A0(net324),
    .A1(net184),
    .A2(net186),
    .A3(net204),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[1] ),
    .A1(\Tile_X0Y0_S4BEG[1] ),
    .A2(net339),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q1 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[322] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0  (.A0(net325),
    .A1(net181),
    .A2(net221),
    .A3(net201),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S4BEG[2] ),
    .A1(\Tile_X0Y0_SS4BEG[2] ),
    .A2(net340),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[326] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0  (.A0(net326),
    .A1(net182),
    .A2(net188),
    .A3(net204),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[3] ),
    .A1(\Tile_X0Y0_S4BEG[3] ),
    .A2(net341),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[330] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0  (.A0(net289),
    .A1(net183),
    .A2(net189),
    .A3(net201),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[4] ),
    .A1(\Tile_X0Y0_S4BEG[0] ),
    .A2(net342),
    .A3(net374),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[334] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net290),
    .A2(net182),
    .A3(net190),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S2BEGb[5] ),
    .A2(net335),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[338] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net291),
    .A2(net183),
    .A3(net191),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[2] ),
    .A1(\Tile_X0Y0_S2BEGb[6] ),
    .A2(net334),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[342] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net292),
    .A2(net184),
    .A3(net192),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[3] ),
    .A1(\Tile_X0Y0_S2BEGb[7] ),
    .A2(net335),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[346] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net285),
    .A2(net181),
    .A3(net185),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S2BEGb[0] ),
    .A2(net334),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(net763),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[350] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net286),
    .A2(net186),
    .A3(net204),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[1] ),
    .A1(\Tile_X0Y0_S4BEG[1] ),
    .A2(net339),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q1 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[354] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net287),
    .A2(net187),
    .A3(net201),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[2] ),
    .A1(\Tile_X0Y0_S4BEG[2] ),
    .A2(net340),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[358] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net288),
    .A2(net188),
    .A3(net204),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[3] ),
    .A1(\Tile_X0Y0_S4BEG[3] ),
    .A2(net341),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[362] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net289),
    .A2(net189),
    .A3(net201),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[4] ),
    .A1(\Tile_X0Y0_S4BEG[0] ),
    .A2(net342),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[366] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net290),
    .A2(net182),
    .A3(net190),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(\Tile_X0Y0_S2BEGb[5] ),
    .A3(net335),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[370] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net291),
    .A2(net183),
    .A3(net191),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(\Tile_X0Y0_S2BEGb[6] ),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[374] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[375] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net292),
    .A2(net184),
    .A3(net192),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(\Tile_X0Y0_S2BEGb[7] ),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[378] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[379] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net285),
    .A2(net181),
    .A3(net185),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(\Tile_X0Y0_S2BEGb[0] ),
    .A3(net334),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(net763),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[382] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[383] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0  (.A0(net184),
    .A1(net337),
    .A2(\Tile_X0Y1_DSP_bot/Q0 ),
    .A3(net764),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/Q3 ),
    .A2(\Tile_X0Y1_DSP_bot/Q4 ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q6 ),
    .A1(\Tile_X0Y1_DSP_bot/Q7 ),
    .A2(\Tile_X0Y1_DSP_bot/Q8 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[112] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net736));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0  (.A0(net183),
    .A1(net336),
    .A2(\Tile_X0Y1_DSP_bot/Q0 ),
    .A3(net764),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/Q3 ),
    .A2(\Tile_X0Y1_DSP_bot/Q4 ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q6 ),
    .A1(\Tile_X0Y1_DSP_bot/Q7 ),
    .A2(\Tile_X0Y1_DSP_bot/Q8 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[116] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net737));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst0  (.A0(net299),
    .A1(net193),
    .A2(net199),
    .A3(\Tile_X0Y0_S2BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst1  (.A0(net346),
    .A1(\Tile_X0Y1_DSP_bot/JN2BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/JS2BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/JW2BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/JW2BEG[5] ),
    .A2(net765),
    .A3(net766),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__conb_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst3_765  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net765));
 sky130_fd_sc_hd__conb_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst3_766  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net766));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[158] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/clr ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_A0  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[0] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[118] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/A0 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_A1  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[120] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/A1 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_A2  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[122] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/A2 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_A3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[124] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/A3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_B0  (.A0(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[0] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[126] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/B0 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_B1  (.A0(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[128] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/B1 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_B2  (.A0(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[130] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/B2 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_B3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[132] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/B3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C0  (.A0(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[0] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[134] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C1  (.A0(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[136] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C2  (.A0(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[138] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C2 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[140] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C4  (.A0(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[0] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[142] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C4 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C5  (.A0(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[144] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C5 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C6  (.A0(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[146] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C6 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C7  (.A0(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[148] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/C7 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_E1BEG0  (.A0(\Tile_X0Y1_DSP_bot/Q3 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[34] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net583));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_E1BEG1  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[36] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_E1BEG2  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[38] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net585));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_E1BEG3  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[40] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0  (.A0(net291),
    .A1(net191),
    .A2(\Tile_X0Y0_SS4BEG[3] ),
    .A3(net344),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[224] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1  (.A0(net317),
    .A1(net187),
    .A2(\Tile_X0Y0_S2BEGb[2] ),
    .A3(net340),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[226] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2  (.A0(net289),
    .A1(net213),
    .A2(\Tile_X0Y0_S2BEGb[4] ),
    .A3(net342),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[228] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3  (.A0(net285),
    .A1(net185),
    .A2(\Tile_X0Y0_S2BEGb[0] ),
    .A3(net375),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[230] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0  (.A0(net326),
    .A1(net191),
    .A2(\Tile_X0Y0_S2BEGb[6] ),
    .A3(net344),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[232] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1  (.A0(net287),
    .A1(net187),
    .A2(\Tile_X0Y0_S2BEGb[2] ),
    .A3(net374),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[234] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2  (.A0(net289),
    .A1(net189),
    .A2(\Tile_X0Y0_SS4BEG[2] ),
    .A3(net342),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[236] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3  (.A0(net285),
    .A1(net220),
    .A2(\Tile_X0Y0_S2BEGb[0] ),
    .A3(net338),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[238] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0  (.A0(net292),
    .A1(net221),
    .A2(\Tile_X0Y0_S2BEGb[7] ),
    .A3(net345),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[240] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1  (.A0(net288),
    .A1(net188),
    .A2(\Tile_X0Y0_S2BEGb[3] ),
    .A3(net373),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[242] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2  (.A0(net290),
    .A1(net190),
    .A2(\Tile_X0Y0_SS4BEG[1] ),
    .A3(net343),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[244] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3  (.A0(net325),
    .A1(net186),
    .A2(\Tile_X0Y0_S2BEGb[1] ),
    .A3(net339),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[246] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0  (.A0(net292),
    .A1(net192),
    .A2(\Tile_X0Y0_S2BEGb[7] ),
    .A3(net366),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[248] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1  (.A0(net288),
    .A1(net188),
    .A2(\Tile_X0Y0_SS4BEG[0] ),
    .A3(net341),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[250] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2  (.A0(net324),
    .A1(net190),
    .A2(\Tile_X0Y0_S2BEGb[5] ),
    .A3(net343),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[252] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3  (.A0(net286),
    .A1(net222),
    .A2(\Tile_X0Y0_S2BEGb[1] ),
    .A3(net339),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[254] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0  (.A0(net299),
    .A1(\Tile_X0Y0_S2BEG[6] ),
    .A2(net352),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[160] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1  (.A0(net195),
    .A1(\Tile_X0Y0_S2BEG[2] ),
    .A2(net348),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[162] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2  (.A0(net297),
    .A1(net197),
    .A2(net350),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[164] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3  (.A0(net293),
    .A1(net193),
    .A2(\Tile_X0Y0_S2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[166] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0  (.A0(net300),
    .A1(net200),
    .A2(\Tile_X0Y0_S2BEG[7] ),
    .A3(net353),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[192] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1  (.A0(net296),
    .A1(net196),
    .A2(\Tile_X0Y0_S2BEG[3] ),
    .A3(net349),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[194] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2  (.A0(net298),
    .A1(net198),
    .A2(\Tile_X0Y0_S2BEG[5] ),
    .A3(net351),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[196] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3  (.A0(net294),
    .A1(net194),
    .A2(\Tile_X0Y0_S2BEG[1] ),
    .A3(net347),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[198] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0  (.A0(net199),
    .A1(\Tile_X0Y0_S2BEG[6] ),
    .A2(net352),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[168] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1  (.A0(net295),
    .A1(net195),
    .A2(net348),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[170] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2  (.A0(net297),
    .A1(net197),
    .A2(\Tile_X0Y0_S2BEG[4] ),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[172] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3  (.A0(net293),
    .A1(\Tile_X0Y0_S2BEG[0] ),
    .A2(net346),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[174] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0  (.A0(net300),
    .A1(net200),
    .A2(\Tile_X0Y0_S2BEG[7] ),
    .A3(net353),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[200] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1  (.A0(net296),
    .A1(net196),
    .A2(\Tile_X0Y0_S2BEG[3] ),
    .A3(net349),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[202] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2  (.A0(net298),
    .A1(net198),
    .A2(\Tile_X0Y0_S2BEG[5] ),
    .A3(net351),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[204] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3  (.A0(net294),
    .A1(net194),
    .A2(\Tile_X0Y0_S2BEG[1] ),
    .A3(net347),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[206] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0  (.A0(net299),
    .A1(net199),
    .A2(net352),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[5] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[176] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1  (.A0(net295),
    .A1(net195),
    .A2(\Tile_X0Y0_S2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[5] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[178] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2  (.A0(net297),
    .A1(\Tile_X0Y0_S2BEG[4] ),
    .A2(net350),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[5] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[180] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3  (.A0(net193),
    .A1(\Tile_X0Y0_S2BEG[0] ),
    .A2(net346),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[5] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[182] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0  (.A0(net300),
    .A1(net200),
    .A2(\Tile_X0Y0_S2BEG[7] ),
    .A3(net353),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[208] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1  (.A0(net296),
    .A1(net196),
    .A2(\Tile_X0Y0_S2BEG[3] ),
    .A3(net349),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[210] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2  (.A0(net298),
    .A1(net198),
    .A2(\Tile_X0Y0_S2BEG[5] ),
    .A3(net351),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[212] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3  (.A0(net294),
    .A1(net194),
    .A2(\Tile_X0Y0_S2BEG[1] ),
    .A3(net347),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[214] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0  (.A0(net299),
    .A1(net199),
    .A2(\Tile_X0Y0_S2BEG[6] ),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[184] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1  (.A0(net295),
    .A1(\Tile_X0Y0_S2BEG[2] ),
    .A2(net348),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[186] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2  (.A0(net197),
    .A1(\Tile_X0Y0_S2BEG[4] ),
    .A2(net350),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[188] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3  (.A0(net293),
    .A1(net193),
    .A2(net346),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[190] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0  (.A0(net300),
    .A1(net200),
    .A2(\Tile_X0Y0_S2BEG[7] ),
    .A3(net353),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[216] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1  (.A0(net296),
    .A1(net196),
    .A2(\Tile_X0Y0_S2BEG[3] ),
    .A3(net349),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[218] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2  (.A0(net298),
    .A1(net198),
    .A2(\Tile_X0Y0_S2BEG[5] ),
    .A3(net351),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[220] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3  (.A0(net294),
    .A1(net194),
    .A2(\Tile_X0Y0_S2BEG[1] ),
    .A3(net347),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[222] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0  (.A0(net326),
    .A1(\Tile_X0Y0_S4BEG[3] ),
    .A2(net366),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[384] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[385] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1  (.A0(net221),
    .A1(\Tile_X0Y0_S4BEG[2] ),
    .A2(net345),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[386] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[387] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2  (.A0(net308),
    .A1(net204),
    .A2(net357),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[388] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[389] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3  (.A0(net301),
    .A1(net201),
    .A2(\Tile_X0Y0_S4BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[390] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[391] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0  (.A0(net188),
    .A1(\Tile_X0Y0_SS4BEG[3] ),
    .A2(net374),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[392] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[393] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1  (.A0(net309),
    .A1(net187),
    .A2(net345),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[394] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[395] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2  (.A0(net324),
    .A1(net220),
    .A2(\Tile_X0Y0_S4BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[396] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[397] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3  (.A0(net301),
    .A1(\Tile_X0Y0_SS4BEG[0] ),
    .A2(net354),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[398] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[399] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0  (.A0(net310),
    .A1(net188),
    .A2(net341),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[400] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[401] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1  (.A0(net325),
    .A1(net187),
    .A2(\Tile_X0Y0_S4BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[402] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[403] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2  (.A0(net308),
    .A1(\Tile_X0Y0_SS4BEG[1] ),
    .A2(net342),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[404] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[405] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3  (.A0(net222),
    .A1(\Tile_X0Y0_S4BEG[0] ),
    .A2(net373),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[406] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[407] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0  (.A0(net310),
    .A1(net213),
    .A2(\Tile_X0Y0_S4BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[408] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[409] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1  (.A0(net309),
    .A1(\Tile_X0Y0_SS4BEG[2] ),
    .A2(net340),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[410] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[411] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2  (.A0(net204),
    .A1(\Tile_X0Y0_S4BEG[1] ),
    .A2(net375),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[412] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[413] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3  (.A0(net317),
    .A1(net201),
    .A2(net338),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[414] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[415] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N1BEG0  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[6] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N1BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N1BEG1  (.A0(\Tile_X0Y1_DSP_bot/Q3 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[8] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N1BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N1BEG2  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[10] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N1BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N1BEG3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[12] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N1BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N4BEG0  (.A0(net287),
    .A1(net308),
    .A2(net204),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[14] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N4BEG1  (.A0(net288),
    .A1(net309),
    .A2(net201),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[16] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N4BEG2  (.A0(net285),
    .A1(net310),
    .A2(net357),
    .A3(net763),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[18] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N4BEG3  (.A0(net286),
    .A1(net301),
    .A2(net354),
    .A3(\Tile_X0Y1_DSP_bot/Q7 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[20] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S1BEG0  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[62] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net663));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S1BEG1  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[64] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net664));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S1BEG2  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[66] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net665));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S1BEG3  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[68] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net666));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S4BEG0  (.A0(net204),
    .A1(\Tile_X0Y0_S2BEGb[2] ),
    .A2(\Tile_X0Y0_S4BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/Q0 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[70] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S4BEG1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[3] ),
    .A2(\Tile_X0Y0_S4BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/Q1 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[72] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net687));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S4BEG2  (.A0(\Tile_X0Y0_S2BEGb[0] ),
    .A1(\Tile_X0Y0_S4BEG[3] ),
    .A2(net357),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[74] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net688));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S4BEG3  (.A0(\Tile_X0Y0_S2BEGb[1] ),
    .A1(\Tile_X0Y0_S4BEG[0] ),
    .A2(net354),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[76] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net689));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_W1BEG0  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[90] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net715));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_W1BEG1  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[92] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net716));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_W1BEG2  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[94] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net717));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_W1BEG3  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[96] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_DSP_bot/JN2BEG[4] ),
    .A1(\Tile_X0Y1_DSP_bot/JN2BEG[6] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[4] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[150] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/JS2BEG[4] ),
    .A1(\Tile_X0Y1_DSP_bot/JS2BEG[6] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[4] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[150] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[152] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/C8 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_DSP_bot/JN2BEG[5] ),
    .A1(\Tile_X0Y1_DSP_bot/JN2BEG[7] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[5] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[7] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[153] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/JS2BEG[5] ),
    .A1(\Tile_X0Y1_DSP_bot/JS2BEG[7] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[5] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[7] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[153] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[155] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/C9 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net183),
    .A2(\Tile_X0Y0_S1BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[42] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[42] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[44] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net618));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net184),
    .A2(\Tile_X0Y0_S1BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[45] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[45] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[47] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net619));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net181),
    .A2(\Tile_X0Y0_S1BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[48] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q8 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[48] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[50] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net620));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net182),
    .A2(\Tile_X0Y0_S1BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[51] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q9 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[51] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[53] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net621));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net183),
    .A2(net336),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[22] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[22] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[24] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_NN4BEG[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net184),
    .A2(net337),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[25] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[25] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[27] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_NN4BEG[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net181),
    .A2(net334),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[28] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q8 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[28] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[30] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_NN4BEG[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net182),
    .A2(net335),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[31] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q9 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[31] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[33] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_NN4BEG[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net183),
    .A2(net336),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[78] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[78] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[80] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net702));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net184),
    .A2(net337),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[81] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[81] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[83] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net703));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net181),
    .A2(net334),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[84] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q8 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[84] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[86] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net704));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net182),
    .A2(net335),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[87] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q9 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[87] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[89] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net705));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0  (.A0(net283),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(net336),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[98] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q6 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[98] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[100] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net750));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0  (.A0(net284),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(net337),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[101] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[101] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[103] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net751));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0  (.A0(net281),
    .A1(\Tile_X0Y0_S1BEG[0] ),
    .A2(net334),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[104] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q8 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[104] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[106] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net752));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0  (.A0(net282),
    .A1(\Tile_X0Y0_S1BEG[1] ),
    .A2(net335),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[107] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q9 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[107] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[109] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net753));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0843_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0844_  (.A0(\Tile_X0Y1_DSP_bot/C0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[0] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0022_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0845_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0022_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[0] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0023_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0846_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0847_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0848_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0849_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[0] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0850_  (.A1(\Tile_X0Y1_DSP_bot/A0 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0851_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0852_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[0] ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0853_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .B_N(\Tile_X0Y1_DSP_bot/B0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0031_ ));
 sky130_fd_sc_hd__nand2_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0854_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0031_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0855_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0856_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0023_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0857_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0023_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0035_ ));
 sky130_fd_sc_hd__or3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0858_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0035_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0036_ ));
 sky130_fd_sc_hd__a21bo_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0859_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[0] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0036_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q0 ));
 sky130_fd_sc_hd__buf_6 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0860_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0861_  (.A(\Tile_X0Y1_DSP_bot/A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0862_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0039_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0863_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0039_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0864_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0865_  (.A(\Tile_X0Y1_DSP_bot/B1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0042_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0866_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0043_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0867_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0042_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0043_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0868_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0869_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0870_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0871_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .A2(\Tile_X0Y1_DSP_bot/B0 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0872_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0039_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0873_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .A2(\Tile_X0Y1_DSP_bot/B1 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0043_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0874_  (.A1(\Tile_X0Y1_DSP_bot/A0 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ));
 sky130_fd_sc_hd__or4_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0875_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0876_  (.A0(\Tile_X0Y1_DSP_bot/C1 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[1] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0053_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0877_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0053_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[1] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0878_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0055_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0879_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0056_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0880_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0055_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0056_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0057_ ));
 sky130_fd_sc_hd__xnor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0881_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0057_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0058_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0882_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0059_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0883_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0058_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0059_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Q1 ));
 sky130_fd_sc_hd__a32o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0884_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0057_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0060_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0885_  (.A(\Tile_X0Y1_DSP_bot/A2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0061_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0886_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0062_ ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0887_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0061_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0062_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ));
 sky130_fd_sc_hd__and2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0888_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ));
 sky130_fd_sc_hd__nor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0889_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0890_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0066_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0891_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0892_  (.A(\Tile_X0Y1_DSP_bot/B2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0068_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0893_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0069_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0894_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0068_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0069_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0895_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0896_  (.A1(\Tile_X0Y1_DSP_bot/A0 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0072_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0897_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0061_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0062_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0898_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0899_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0900_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ));
 sky130_fd_sc_hd__o311a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0901_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0066_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0072_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0077_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0902_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0078_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0903_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ));
 sky130_fd_sc_hd__o21a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0904_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0068_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0069_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ));
 sky130_fd_sc_hd__o2bb2a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0905_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0078_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0081_ ));
 sky130_fd_sc_hd__nor3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0906_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0077_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0081_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0907_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0077_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0081_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0083_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0908_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0083_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0084_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0909_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0910_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0911_  (.A0(\Tile_X0Y1_DSP_bot/C2 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[2] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0087_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0912_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[2] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0088_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0913_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0087_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0088_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0089_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0914_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0084_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0089_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0090_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0915_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0084_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0089_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0091_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0916_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0090_ ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0091_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0092_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0917_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0060_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0092_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0093_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0918_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0919_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0093_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[2] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0095_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0920_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0095_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q2 ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0921_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[3] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0096_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0922_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .A2(\Tile_X0Y1_DSP_bot/C3 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0096_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0097_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0923_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0098_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0924_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0097_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0098_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0099_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0925_  (.A(\Tile_X0Y1_DSP_bot/B3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0100_ ));
 sky130_fd_sc_hd__nand2_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0926_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0927_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0100_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0928_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0929_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0104_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0930_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0072_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0104_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0066_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ));
 sky130_fd_sc_hd__buf_6 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0931_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0932_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0933_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/A3 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0934_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0935_  (.A(\Tile_X0Y1_DSP_bot/A3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0110_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0936_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0111_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0937_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0110_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0111_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ));
 sky130_fd_sc_hd__buf_6 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0938_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0939_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ));
 sky130_fd_sc_hd__o2111ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0940_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0115_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0941_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0116_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0942_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0115_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0116_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0943_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0118_ ));
 sky130_fd_sc_hd__a22oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0944_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0119_ ));
 sky130_fd_sc_hd__o21bai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0945_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0118_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0119_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0120_ ));
 sky130_fd_sc_hd__nand4_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0946_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0120_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0947_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0120_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0948_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0949_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ));
 sky130_fd_sc_hd__or3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0950_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0099_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0951_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0099_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0126_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0952_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0060_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0091_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0090_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0953_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0126_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0128_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0954_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0126_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0129_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0955_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0128_ ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0129_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0130_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0956_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0130_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[3] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0131_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0957_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0131_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q3 ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0958_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B_N(\Tile_X0Y1_DSP_bot/B3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0959_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0133_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0960_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0115_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0116_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0134_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0961_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0133_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0134_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0962_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0963_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/A4 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0964_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0965_  (.A(\Tile_X0Y1_DSP_bot/A4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0139_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0966_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0140_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0967_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0139_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0140_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ));
 sky130_fd_sc_hd__nor2b_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0968_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B_N(\Tile_X0Y1_DSP_bot/B2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ));
 sky130_fd_sc_hd__and2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0969_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0970_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0144_ ));
 sky130_fd_sc_hd__a41oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0971_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0144_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0972_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0973_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0974_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0148_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0975_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0976_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0150_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0977_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .B(\Tile_X0Y1_DSP_bot/B4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0978_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[4] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ));
 sky130_fd_sc_hd__a32o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0979_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0153_ ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0980_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0100_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0981_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/B4 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ));
 sky130_fd_sc_hd__or4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0982_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0156_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0983_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0156_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ));
 sky130_fd_sc_hd__a221o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0984_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0985_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0148_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0150_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0153_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0986_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0160_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0987_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0161_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0988_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0162_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0989_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0161_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0162_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0150_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0990_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0153_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0991_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0160_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0992_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0993_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0167_ ));
 sky130_fd_sc_hd__a32o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0994_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0167_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0168_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0995_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0169_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0996_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0170_ ));
 sky130_fd_sc_hd__a311o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0997_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0169_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0170_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0998_  (.A0(\Tile_X0Y1_DSP_bot/C4 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[4] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0172_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0999_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0172_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[4] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0173_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1000_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0168_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0174_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1001_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0174_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0175_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1002_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0168_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ));
 sky130_fd_sc_hd__o221a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1003_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0097_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0098_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0177_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1004_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0177_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1005_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0175_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0179_ ));
 sky130_fd_sc_hd__or3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1006_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0175_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0180_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1007_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0179_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0180_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0181_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1008_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0181_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[4] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0182_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1009_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0182_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q4 ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1010_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0174_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0183_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1011_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ));
 sky130_fd_sc_hd__and4_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1012_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0167_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1013_  (.A(\Tile_X0Y1_DSP_bot/A5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0186_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1014_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0187_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1015_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0186_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1016_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ));
 sky130_fd_sc_hd__a41oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1017_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1018_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1019_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ),
    .A2(\Tile_X0Y1_DSP_bot/A5 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1020_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1021_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1022_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1023_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .B(\Tile_X0Y1_DSP_bot/A3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1024_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1025_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1026_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1027_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0200_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1028_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0201_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1029_  (.A(\Tile_X0Y1_DSP_bot/B4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0202_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1030_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0203_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1031_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0202_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0203_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1032_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1033_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1034_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ));
 sky130_fd_sc_hd__or2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1035_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[5] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1036_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B5 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0209_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1037_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0209_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0210_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1038_  (.A(\Tile_X0Y1_DSP_bot/B5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0211_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1039_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0212_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1040_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0211_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0212_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1041_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1042_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1043_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0210_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1044_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0200_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0201_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1045_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0218_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1046_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0219_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1047_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0218_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0219_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0200_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0220_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1048_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0220_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1049_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ));
 sky130_fd_sc_hd__o211a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1050_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1051_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0224_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1052_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0225_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1053_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0224_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0225_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1054_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1055_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ));
 sky130_fd_sc_hd__o22a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1056_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0229_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1057_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1058_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ));
 sky130_fd_sc_hd__a41o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1059_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0232_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1060_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0229_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0232_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0219_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0233_ ));
 sky130_fd_sc_hd__o41a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1061_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0234_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1062_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0233_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0234_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1063_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0236_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1064_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0236_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0237_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1065_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0237_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1066_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1067_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0240_ ));
 sky130_fd_sc_hd__o2111ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1068_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0241_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1069_  (.A0(\Tile_X0Y1_DSP_bot/C5 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[5] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0242_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1070_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0242_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[5] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0243_ ));
 sky130_fd_sc_hd__a21boi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1071_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0240_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0241_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0243_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0244_ ));
 sky130_fd_sc_hd__and3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1072_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0243_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0241_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0240_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0245_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1073_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0244_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0245_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0246_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1074_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0183_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0246_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0247_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1075_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0247_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[5] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0248_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1076_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0248_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q5 ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1077_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0183_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0245_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0244_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0249_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1078_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0224_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0225_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1079_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0251_ ));
 sky130_fd_sc_hd__a2111o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1080_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0251_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0169_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0170_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0252_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1081_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0253_ ));
 sky130_fd_sc_hd__o211ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1082_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0254_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1083_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0229_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1084_  (.A(\Tile_X0Y1_DSP_bot/A6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0256_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1085_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0257_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1086_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0256_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0257_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1087_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1088_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0260_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1089_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0260_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1090_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/A5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0262_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1091_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0262_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1092_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0264_ ));
 sky130_fd_sc_hd__nor2b_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1093_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B_N(\Tile_X0Y1_DSP_bot/A6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1094_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0266_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1095_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0266_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1096_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0031_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ));
 sky130_fd_sc_hd__and2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1097_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ));
 sky130_fd_sc_hd__nor2b_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1098_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B_N(\Tile_X0Y1_DSP_bot/A4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1099_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1100_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0264_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1101_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ),
    .A2(\Tile_X0Y1_DSP_bot/A6 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0257_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1102_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1103_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1104_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0276_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1105_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0264_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0277_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1106_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0278_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1107_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B2 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0279_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1108_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0278_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0279_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0280_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1109_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0277_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0280_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0281_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1110_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1111_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ));
 sky130_fd_sc_hd__a22o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1112_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1113_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ));
 sky130_fd_sc_hd__o2111a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1114_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0276_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0281_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1115_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0287_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1116_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0287_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0288_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1117_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0277_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0280_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1118_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1119_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0288_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1120_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1121_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[6] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ));
 sky130_fd_sc_hd__o21a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1122_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/B6 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1123_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1124_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0296_ ));
 sky130_fd_sc_hd__a31oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1125_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0296_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1126_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1127_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B6 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1128_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ));
 sky130_fd_sc_hd__o2bb2a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1129_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1130_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0288_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0302_ ));
 sky130_fd_sc_hd__o22a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1131_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0220_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1132_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0302_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1133_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1134_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0276_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0281_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ));
 sky130_fd_sc_hd__o211a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1135_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1136_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0308_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1137_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0308_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1138_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0310_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1139_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0311_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1140_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0310_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0311_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0312_ ));
 sky130_fd_sc_hd__o21bai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1141_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0312_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1142_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0237_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0251_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0314_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1143_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0314_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0315_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1144_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0254_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0315_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0316_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1145_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0317_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1146_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0317_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1147_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ));
 sky130_fd_sc_hd__a221oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1148_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0310_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0311_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0317_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0320_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1149_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1150_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0312_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0322_ ));
 sky130_fd_sc_hd__o21bai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1151_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0320_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0322_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0314_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0323_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1152_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0323_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0324_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1153_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0252_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0253_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0316_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0324_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1154_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0326_ ));
 sky130_fd_sc_hd__nor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1155_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1156_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0328_ ));
 sky130_fd_sc_hd__a2bb2oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1157_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0328_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0329_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1158_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0329_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0315_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0330_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1159_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0326_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0330_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1160_  (.A0(\Tile_X0Y1_DSP_bot/C6 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[6] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0332_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1161_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0332_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0333_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1162_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[6] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0334_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1163_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0333_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0334_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0335_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1164_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0333_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0334_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0336_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1165_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0336_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0337_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1166_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0335_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0337_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0338_ ));
 sky130_fd_sc_hd__xor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1167_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0249_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0338_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0339_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1168_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0340_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1169_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0339_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0340_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Q6 ));
 sky130_fd_sc_hd__a32oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1170_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0336_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0249_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0335_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1171_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0326_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0330_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1172_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B5 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1173_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0344_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1174_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0344_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ));
 sky130_fd_sc_hd__or2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1175_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[7] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ));
 sky130_fd_sc_hd__o21a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1176_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B7 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1177_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1178_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ));
 sky130_fd_sc_hd__and4b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1179_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0350_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1180_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B7 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1181_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0352_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1182_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0352_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1183_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0354_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1184_  (.A(\Tile_X0Y1_DSP_bot/A7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0355_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1185_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0356_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1186_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0355_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0356_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1187_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1188_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ),
    .A2(\Tile_X0Y1_DSP_bot/A7 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0356_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1189_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1190_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0361_ ));
 sky130_fd_sc_hd__o2111a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1191_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0362_ ));
 sky130_fd_sc_hd__a22oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1192_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0363_ ));
 sky130_fd_sc_hd__o32a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1193_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0363_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0364_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1194_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0361_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0362_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0364_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1195_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ));
 sky130_fd_sc_hd__a41o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1196_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0367_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1197_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1198_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0363_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1199_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1200_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0367_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1201_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1202_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B5 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0373_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1203_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0374_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1204_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0374_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ));
 sky130_fd_sc_hd__a22oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1205_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0376_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1206_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0373_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0376_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1207_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1208_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1209_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ));
 sky130_fd_sc_hd__a41o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1210_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ));
 sky130_fd_sc_hd__o22a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1211_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1212_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ));
 sky130_fd_sc_hd__o2111ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1213_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0384_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1214_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0385_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1215_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0287_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0386_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1216_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0385_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0386_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1217_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0384_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0388_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1218_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1219_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0367_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1220_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1221_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0350_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0354_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0388_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0392_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1222_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0393_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1223_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0394_ ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1224_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0393_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0394_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1225_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1226_  (.A1(\Tile_X0Y1_DSP_bot/A0 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1227_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1228_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0399_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1229_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0400_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1230_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0392_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0399_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0400_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0401_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1231_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0402_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1232_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0403_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1233_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0402_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0403_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0404_ ));
 sky130_fd_sc_hd__o22a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1234_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0385_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0386_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0405_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1235_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0406_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1236_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0404_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0405_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0406_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1237_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0408_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1238_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0408_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1239_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ));
 sky130_fd_sc_hd__o32ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1240_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0401_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1241_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0412_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1242_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0406_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0412_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0413_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1243_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0400_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0392_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0399_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ));
 sky130_fd_sc_hd__a211oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1244_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1245_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0413_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1246_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0329_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ));
 sky130_fd_sc_hd__o221a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1247_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0418_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1248_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0418_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0419_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1249_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0419_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0420_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1250_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0420_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0421_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1251_  (.A0(\Tile_X0Y1_DSP_bot/C7 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[7] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0422_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1252_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1253_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0422_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[7] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1254_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0421_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0425_ ));
 sky130_fd_sc_hd__xor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1255_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0425_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0426_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1256_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0426_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[7] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0427_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1257_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0427_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q7 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1258_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ));
 sky130_fd_sc_hd__or3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1259_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0429_ ));
 sky130_fd_sc_hd__o311a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1260_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0405_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0393_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0394_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0430_ ));
 sky130_fd_sc_hd__o22a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1261_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0431_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1262_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0430_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0431_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0432_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1263_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0432_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0433_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1264_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0429_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0433_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0434_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1265_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0434_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ));
 sky130_fd_sc_hd__o32ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1266_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0431_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0430_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0429_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0401_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0436_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1267_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0437_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1268_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1269_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1270_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1271_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0441_ ));
 sky130_fd_sc_hd__o32ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1272_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0441_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ));
 sky130_fd_sc_hd__o211a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1273_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1274_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1275_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ));
 sky130_fd_sc_hd__a41oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1276_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1277_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .B_N(\Tile_X0Y1_DSP_bot/B4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0447_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1278_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0203_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0447_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1279_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ));
 sky130_fd_sc_hd__nand2_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1280_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1281_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1282_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ));
 sky130_fd_sc_hd__a32o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1283_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1284_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ));
 sky130_fd_sc_hd__nand2_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1285_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1286_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0456_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1287_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0456_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1288_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0458_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1289_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0459_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1290_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0459_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0362_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1291_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0458_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1292_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0462_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1293_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0462_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1294_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1295_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0465_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1296_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1297_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0465_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1298_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0468_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1299_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0469_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1300_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0374_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0469_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0470_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1301_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B6 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0471_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1302_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0468_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0470_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0471_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1303_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1304_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0474_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1305_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0475_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1306_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0474_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0475_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1307_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0477_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1308_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B7 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1309_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0479_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1310_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0480_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1311_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0481_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1312_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0479_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0480_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0481_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0482_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1313_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0437_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0477_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0482_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1314_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0458_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1315_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0462_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0485_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1316_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0486_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1317_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0485_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0486_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0487_ ));
 sky130_fd_sc_hd__a21o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1318_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0487_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1319_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0474_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0475_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0489_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1320_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0489_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ));
 sky130_fd_sc_hd__a31o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1321_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ));
 sky130_fd_sc_hd__a21o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1322_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1323_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1324_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0436_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ));
 sky130_fd_sc_hd__a221o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1325_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0432_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0495_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1326_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0495_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1327_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0495_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1328_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1329_  (.A0(\Tile_X0Y1_DSP_bot/C8 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[8] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0499_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1330_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[8] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0500_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1331_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0499_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0500_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1332_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0502_ ));
 sky130_fd_sc_hd__or3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1333_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0503_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1334_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0502_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0503_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0504_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1335_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0413_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0505_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1336_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0505_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0506_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1337_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0506_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0507_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1338_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0420_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0507_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0508_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1339_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0421_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0509_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1340_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0508_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0509_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0510_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1341_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0504_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0510_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0511_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1342_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0510_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0504_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0512_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1343_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0513_ ));
 sky130_fd_sc_hd__a31o_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1344_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0511_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0512_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0513_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q8 ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1345_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0508_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0509_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0514_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1346_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0515_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1347_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0514_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0502_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0515_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ));
 sky130_fd_sc_hd__a32oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1348_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0505_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0517_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1349_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0436_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0518_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1350_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0517_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0518_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1351_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0520_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1352_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1353_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0522_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1354_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ));
 sky130_fd_sc_hd__nand4_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1355_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0524_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1356_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .A2(\Tile_X0Y1_DSP_bot/A4 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1357_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0524_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0526_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1358_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1359_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0528_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1360_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0522_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0526_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0528_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1361_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0524_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0530_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1362_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0531_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1363_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0441_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0532_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1364_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0530_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0531_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0532_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1365_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ));
 sky130_fd_sc_hd__o22a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1366_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0522_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0526_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0528_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1367_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ));
 sky130_fd_sc_hd__a211o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1368_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0537_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1369_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0530_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0531_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0538_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1370_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0537_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0538_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1371_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0540_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1372_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0541_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1373_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0542_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1374_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0540_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0541_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0542_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1375_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0544_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1376_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0544_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1377_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0546_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1378_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0547_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1379_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0546_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0547_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0548_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1380_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0548_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1381_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0550_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1382_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0550_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0551_ ));
 sky130_fd_sc_hd__o2bb2a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1383_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1384_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B7 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0553_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1385_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0553_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ));
 sky130_fd_sc_hd__nor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1386_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0555_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1387_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0551_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0555_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0556_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1388_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0556_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1389_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0487_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0558_ ));
 sky130_fd_sc_hd__a221o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1390_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0559_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1391_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0555_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0559_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1392_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0551_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1393_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0558_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1394_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1395_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1396_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0565_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1397_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0565_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0566_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1398_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0479_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0480_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0567_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1399_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0567_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0481_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0568_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1400_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0568_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1401_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0558_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1402_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0571_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1403_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0572_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1404_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0571_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0572_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1405_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0566_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0574_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1406_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0520_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0574_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0575_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1407_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0520_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0574_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0576_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1408_  (.A0(\Tile_X0Y1_DSP_bot/C9 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[9] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0577_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1409_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0577_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[9] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0578_ ));
 sky130_fd_sc_hd__o21bai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1410_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0575_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0576_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0578_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1411_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0575_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0576_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0580_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1412_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0580_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0578_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1413_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0582_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1414_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0583_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1415_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0582_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0583_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0584_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1416_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0584_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[9] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0585_ ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1417_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0585_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q9 ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1418_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0566_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1419_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0587_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1420_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0588_ ));
 sky130_fd_sc_hd__nand3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1421_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0589_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1422_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0588_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0589_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0590_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1423_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0572_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0590_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1424_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0592_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1425_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0593_ ));
 sky130_fd_sc_hd__a221o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1426_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0593_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1427_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0595_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1428_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .A2(\Tile_X0Y1_DSP_bot/A4 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0595_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1429_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1430_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1431_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1432_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0600_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1433_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0600_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0601_ ));
 sky130_fd_sc_hd__o2111ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1434_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0600_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0602_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1435_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0601_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0602_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1436_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ));
 sky130_fd_sc_hd__or4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1437_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0605_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1438_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0605_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0606_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1439_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0606_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1440_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0608_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1441_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0605_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1442_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0608_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1443_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1444_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ));
 sky130_fd_sc_hd__a21boi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1445_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0553_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1446_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1447_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0559_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0615_ ));
 sky130_fd_sc_hd__a41oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1448_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0556_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0615_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0616_ ));
 sky130_fd_sc_hd__nand3b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1449_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0617_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1450_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0616_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0617_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0618_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1451_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0619_ ));
 sky130_fd_sc_hd__nor3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1452_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0619_ ),
    .C_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0620_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1453_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0621_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1454_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0620_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0621_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0622_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1455_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0618_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0622_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1456_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0587_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0592_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ));
 sky130_fd_sc_hd__a32oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1457_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1458_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1459_  (.A0(\Tile_X0Y1_DSP_bot/C10 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[10] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0627_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1460_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0627_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0628_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1461_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[10] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0629_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1462_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0628_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0629_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0630_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1463_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0628_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0629_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0631_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1464_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0631_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1465_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0630_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0633_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1466_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0633_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1467_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0635_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1468_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0630_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0635_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0636_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1469_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0637_ ));
 sky130_fd_sc_hd__a31o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1470_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0636_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0637_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q10 ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1471_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0631_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0638_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1472_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0633_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1473_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0640_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1474_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0616_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0617_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0640_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1475_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0642_ ));
 sky130_fd_sc_hd__a31o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1476_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0643_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1477_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0209_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0644_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1478_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0645_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1479_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1480_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B(\Tile_X0Y1_DSP_bot/A7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0647_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1481_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0648_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1482_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0647_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0648_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0649_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1483_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0650_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1484_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0649_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0650_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0651_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1485_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0651_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0652_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1486_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0653_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1487_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0649_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0650_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0654_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1488_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0655_ ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1489_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0653_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0654_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0655_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1490_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0652_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1491_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0652_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ));
 sky130_fd_sc_hd__o211ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1492_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0644_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0645_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0659_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1493_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ));
 sky130_fd_sc_hd__a32o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1494_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0661_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1495_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0661_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0662_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1496_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0643_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0659_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0662_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1497_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0644_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0645_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ));
 sky130_fd_sc_hd__a22oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1498_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0661_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0665_ ));
 sky130_fd_sc_hd__a31oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1499_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0666_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1500_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0665_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0666_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1501_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0668_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1502_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0668_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ));
 sky130_fd_sc_hd__a21boi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1503_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1504_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0619_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ));
 sky130_fd_sc_hd__nand3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1505_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1506_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1507_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0674_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1508_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0674_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0675_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1509_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0675_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0676_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1510_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0642_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0676_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1511_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0676_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0678_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1512_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0618_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0678_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1513_  (.A0(\Tile_X0Y1_DSP_bot/C11 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[11] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0680_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1514_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1515_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0680_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[11] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1516_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1517_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0684_ ));
 sky130_fd_sc_hd__nor4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1518_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0638_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0684_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0685_ ));
 sky130_fd_sc_hd__o22a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1519_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0638_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0684_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0686_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1520_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0685_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0686_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0687_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1521_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0687_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[11] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0688_ ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1522_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0688_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q11 ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1523_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0689_ ));
 sky130_fd_sc_hd__a31oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1524_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0689_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0690_ ));
 sky130_fd_sc_hd__o2111a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1525_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0675_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0622_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0691_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1526_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0691_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1527_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0674_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0693_ ));
 sky130_fd_sc_hd__o22ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1528_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0693_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0694_ ));
 sky130_fd_sc_hd__a31oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1529_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0691_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0694_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ));
 sky130_fd_sc_hd__or2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1530_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1531_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1532_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0698_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1533_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1534_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0698_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0700_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1535_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0698_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1536_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0700_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1537_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0700_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0703_ ));
 sky130_fd_sc_hd__o311a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1538_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0655_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0651_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0704_ ));
 sky130_fd_sc_hd__o31a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1539_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0704_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0705_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1540_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0703_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0705_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0706_ ));
 sky130_fd_sc_hd__nor3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1541_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0705_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0703_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1542_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0665_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0666_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0708_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1543_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0708_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0709_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1544_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0706_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0709_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0710_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1545_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0709_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0706_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1546_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0712_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1547_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0710_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0712_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1548_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1549_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0715_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1550_  (.A0(\Tile_X0Y1_DSP_bot/C12 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[12] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0716_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1551_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0716_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0717_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1552_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[12] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0718_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1553_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0717_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0718_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0719_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1554_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0715_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0719_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0720_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1555_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0715_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0719_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0721_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1556_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0720_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0721_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0722_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1557_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0690_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0722_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0723_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1558_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0723_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[12] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0724_ ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1559_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0724_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q12 ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1560_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1561_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0726_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1562_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0727_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1563_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0726_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0727_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ));
 sky130_fd_sc_hd__xor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1564_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0729_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1565_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0729_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1566_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0731_ ));
 sky130_fd_sc_hd__a311o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1567_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0731_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0729_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0732_ ));
 sky130_fd_sc_hd__a211oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1568_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0732_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1569_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0732_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1570_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0735_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1571_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0735_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0736_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1572_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0712_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0737_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1573_  (.A0(\Tile_X0Y1_DSP_bot/C13 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[13] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0738_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1574_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0738_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0739_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1575_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[13] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0740_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1576_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0736_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0737_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0739_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0740_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1577_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0739_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0740_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0742_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1578_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0736_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0737_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0742_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0743_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1579_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0743_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0744_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1580_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0690_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0721_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0720_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0745_ ));
 sky130_fd_sc_hd__xor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1581_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0744_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0745_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0746_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1582_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0746_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[13] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0747_ ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1583_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0747_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q13 ));
 sky130_fd_sc_hd__a211o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1584_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0748_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1585_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0749_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1586_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0748_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0749_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0750_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1587_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0748_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0749_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0751_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1588_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0752_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1589_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0752_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0753_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1590_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0754_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1591_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0750_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0751_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0753_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0754_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1592_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0756_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1593_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0757_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1594_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0756_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0757_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0758_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1595_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0750_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0751_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0759_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1596_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0752_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0758_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0759_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1597_  (.A0(\Tile_X0Y1_DSP_bot/C14 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[14] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0761_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1598_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0761_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[14] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1599_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1600_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1601_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1602_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0766_ ));
 sky130_fd_sc_hd__o41ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1603_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0766_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0717_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0718_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0743_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0767_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1604_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0689_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0768_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1605_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0722_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0769_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1606_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0768_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0769_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0744_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0770_ ));
 sky130_fd_sc_hd__a21boi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1607_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0767_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0770_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1608_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0772_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1609_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0773_ ));
 sky130_fd_sc_hd__a2bb2o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1610_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0772_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0773_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[14] ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q14 ));
 sky130_fd_sc_hd__o221a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1611_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0774_ ));
 sky130_fd_sc_hd__o31ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1612_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0774_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1613_  (.A0(\Tile_X0Y1_DSP_bot/C15 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[15] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0776_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1614_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0776_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[15] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1615_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1616_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0779_ ));
 sky130_fd_sc_hd__o311ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1617_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0774_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0779_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1618_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0781_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1619_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0782_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1620_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0783_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1621_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0782_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0783_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0784_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1622_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0781_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0784_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0785_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1623_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0786_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1624_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0785_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0786_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Q15 ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1625_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1626_  (.A0(\Tile_X0Y1_DSP_bot/C16 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[16] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0788_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1627_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0788_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[16] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0789_ ));
 sky130_fd_sc_hd__xnor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1628_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0789_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1629_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0767_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0791_ ));
 sky130_fd_sc_hd__a32oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1630_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0792_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1631_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0791_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0792_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0793_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1632_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0794_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1633_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0793_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0794_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0770_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1634_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0796_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1635_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0797_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1636_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[16] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0796_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0797_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q16 ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1637_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0789_ ),
    .C(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1638_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1639_  (.A0(\Tile_X0Y1_DSP_bot/C17 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[17] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0800_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1640_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0800_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0801_ ));
 sky130_fd_sc_hd__a221o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1641_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B2(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0801_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1642_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0801_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0803_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1643_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0803_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0804_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1644_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0804_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0805_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1645_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0804_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0806_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1646_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0805_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0806_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0807_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1647_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0807_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q17 ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1648_  (.A0(\Tile_X0Y1_DSP_bot/C18 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[18] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0808_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1649_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0808_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[18] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1650_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1651_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .A2(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0811_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1652_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0812_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1653_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1654_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0803_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ));
 sky130_fd_sc_hd__a22oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1655_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0811_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0812_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1656_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .A2(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0816_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1657_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ),
    .C(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0817_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1658_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0816_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0817_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0818_ ));
 sky130_fd_sc_hd__a31o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1659_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0818_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0819_ ));
 sky130_fd_sc_hd__a2bb2o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1660_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0819_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Q18 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1661_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0820_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1662_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ),
    .C(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0821_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1663_  (.A0(\Tile_X0Y1_DSP_bot/C19 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[19] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0822_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1664_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0822_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[19] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0823_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1665_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0823_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0824_ ));
 sky130_fd_sc_hd__o21bai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1666_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0821_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0824_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0825_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1667_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0817_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0816_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0826_ ));
 sky130_fd_sc_hd__o211ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1668_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0824_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0826_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0827_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1669_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0825_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0827_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0828_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1670_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0820_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0828_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Q19 ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1671_  (.A(\Tile_X0Y1_DSP_bot/clr ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1672_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0035_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0000_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1673_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0058_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0001_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1674_  (.A(\Tile_X0Y1_DSP_bot/clr ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1675_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0093_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0831_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1676_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0831_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0002_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1677_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0130_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0832_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1678_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0832_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0003_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1679_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0833_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1680_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0833_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0004_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1681_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0247_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0834_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1682_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0834_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0005_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1683_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0339_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0006_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1684_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0426_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0835_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1685_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0835_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0007_ ));
 sky130_fd_sc_hd__and3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1686_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0511_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0512_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0836_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1687_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0836_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0008_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1688_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0584_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0837_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1689_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0837_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0009_ ));
 sky130_fd_sc_hd__and3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1690_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0636_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0838_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1691_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0838_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0010_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1692_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0687_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0839_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1693_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0839_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0011_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1694_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0723_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0840_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1695_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0840_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0012_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1696_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0746_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0841_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1697_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0841_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0013_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1698_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0783_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0773_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0014_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1699_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0785_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0015_ ));
 sky130_fd_sc_hd__and3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1700_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0796_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0842_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1701_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0842_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0016_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1702_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0805_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0806_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0017_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1703_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0818_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0020_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1704_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0020_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0018_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1705_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0825_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0827_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0019_ ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1706_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0000_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1707_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0001_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1708_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0002_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1709_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1710_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0004_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[4] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1711_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[5] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1712_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0006_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[6] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1713_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0007_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[7] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1714_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0008_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[8] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1715_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0009_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[9] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1716_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0010_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[10] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1717_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0011_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[11] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1718_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0012_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[12] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1719_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0013_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[13] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1720_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0014_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[14] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1721_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0015_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[15] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1722_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0016_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[16] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1723_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0017_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1724_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0018_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[18] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1725_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0019_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[19] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1726_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1727_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1728_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1729_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1730_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1731_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1732_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1733_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1734_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1735_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1736_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1737_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1738_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1739_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1740_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1741_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1742_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1743_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1744_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1745_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1746_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1747_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1748_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1749_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1750_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1751_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1752_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1753_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1754_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1755_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1756_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1757_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1758_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1759_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1760_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1761_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[19] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[11] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_N4BEG[9] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_0/_0_  (.A(net311),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[0] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_1/_0_  (.A(net312),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_10/_0_  (.A(net306),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_11/_0_  (.A(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_2/_0_  (.A(net313),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/N4END_inbuf_3/_0_  (.A(net314),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[3] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_4/_0_  (.A(net315),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_5/_0_  (.A(net316),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_6/_0_  (.A(net302),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_7/_0_  (.A(net303),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_8/_0_  (.A(net304),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_9/_0_  (.A(net305),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[9] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[11] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[2] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_NN4BEG[9] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_0/_0_  (.A(net327),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_1/_0_  (.A(net328),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/NN4END_inbuf_10/_0_  (.A(net322),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_11/_0_  (.A(net323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[11] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_2/_0_  (.A(net329),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[2] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_3/_0_  (.A(net330),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_4/_0_  (.A(net331),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_5/_0_  (.A(net332),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_6/_0_  (.A(net318),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[6] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_7/_0_  (.A(net319),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_8/_0_  (.A(net320),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_9/_0_  (.A(net321),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_0/_0_  (.A(\Tile_X0Y0_S4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/S4END_inbuf_1/_0_  (.A(\Tile_X0Y0_S4BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/S4END_inbuf_10/_0_  (.A(\Tile_X0Y0_S4BEG[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_11/_0_  (.A(\Tile_X0Y0_S4BEG[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_2/_0_  (.A(\Tile_X0Y0_S4BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_3/_0_  (.A(\Tile_X0Y0_S4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_4/_0_  (.A(\Tile_X0Y0_S4BEG[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_5/_0_  (.A(\Tile_X0Y0_S4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_6/_0_  (.A(\Tile_X0Y0_S4BEG[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[6] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/S4END_inbuf_7/_0_  (.A(\Tile_X0Y0_S4BEG[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[7] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_8/_0_  (.A(\Tile_X0Y0_S4BEG[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[8] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_9/_0_  (.A(\Tile_X0Y0_S4BEG[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_0/_0_  (.A(\Tile_X0Y0_SS4BEG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_1/_0_  (.A(\Tile_X0Y0_SS4BEG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[1] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_10/_0_  (.A(\Tile_X0Y0_SS4BEG[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[10] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/SS4END_inbuf_11/_0_  (.A(\Tile_X0Y0_SS4BEG[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_2/_0_  (.A(\Tile_X0Y0_SS4BEG[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_3/_0_  (.A(\Tile_X0Y0_SS4BEG[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_4/_0_  (.A(\Tile_X0Y0_SS4BEG[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_5/_0_  (.A(\Tile_X0Y0_SS4BEG[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_6/_0_  (.A(\Tile_X0Y0_SS4BEG[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_7/_0_  (.A(\Tile_X0Y0_SS4BEG[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/SS4END_inbuf_8/_0_  (.A(\Tile_X0Y0_SS4BEG[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/SS4END_inbuf_9/_0_  (.A(\Tile_X0Y0_SS4BEG[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_0/_0_  (.A(net358),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_1/_0_  (.A(net359),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_2/_0_  (.A(net360),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_3/_0_  (.A(net361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_4/_0_  (.A(net362),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_5/_0_  (.A(net363),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_6/_0_  (.A(net364),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_7/_0_  (.A(net365),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_8/_0_  (.A(net355),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_9/_0_  (.A(net356),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_0/_0_  (.A(net376),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_1/_0_  (.A(net377),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_10/_0_  (.A(net371),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_11/_0_  (.A(net372),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_2/_0_  (.A(net378),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_3/_0_  (.A(net379),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_4/_0_  (.A(net380),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_5/_0_  (.A(net381),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_6/_0_  (.A(net367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_7/_0_  (.A(net368),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_8/_0_  (.A(net369),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_9/_0_  (.A(net370),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_0/_0_  (.A(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_1/_0_  (.A(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_10/_0_  (.A(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_11/_0_  (.A(net231),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_12/_0_  (.A(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[12] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/data_inbuf_13/_0_  (.A(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_14/_0_  (.A(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_15/_0_  (.A(net235),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_16/_0_  (.A(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_17/_0_  (.A(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_18/_0_  (.A(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_19/_0_  (.A(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_2/_0_  (.A(net251),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_20/_0_  (.A(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[20] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_21/_0_  (.A(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[21] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_22/_0_  (.A(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[22] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_23/_0_  (.A(net244),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[23] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_24/_0_  (.A(net245),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[24] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_25/_0_  (.A(net246),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[25] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_26/_0_  (.A(net247),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[26] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_27/_0_  (.A(net248),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[27] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_28/_0_  (.A(net249),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[28] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_29/_0_  (.A(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[29] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_3/_0_  (.A(net254),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_30/_0_  (.A(net252),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[30] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_31/_0_  (.A(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[31] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_4/_0_  (.A(net255),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_5/_0_  (.A(net256),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_6/_0_  (.A(net257),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_7/_0_  (.A(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_8/_0_  (.A(net259),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_9/_0_  (.A(net260),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_12/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_13/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_14/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_15/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_16/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_17/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_18/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_19/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_20/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_21/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_22/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_23/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_24/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_25/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_26/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_27/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_28/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_29/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_30/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_31/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/inst_clk_buf  (.A(net333),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_UserCLKo));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_0/_0_  (.A(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_1/_0_  (.A(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_10/_0_  (.A(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_11/_0_  (.A(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_12/_0_  (.A(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_13/_0_  (.A(net265),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_14/_0_  (.A(net266),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_15/_0_  (.A(net267),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_16/_0_  (.A(net268),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_17/_0_  (.A(net269),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_18/_0_  (.A(net270),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_19/_0_  (.A(net271),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_2/_0_  (.A(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[2] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_3/_0_  (.A(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_4/_0_  (.A(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_5/_0_  (.A(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_6/_0_  (.A(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_7/_0_  (.A(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[7] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_8/_0_  (.A(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_9/_0_  (.A(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[9] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[0] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[1] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[10] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[11] ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_12/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[12] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/strobe_outbuf_13/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[13] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_14/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[14] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_15/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[15] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_16/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_17/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[17] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_18/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[18] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_19/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[19] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[2] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[3] ));
 sky130_fd_sc_hd__clkbuf_16 \Tile_X0Y1_DSP_bot/strobe_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[4] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[5] ));
 sky130_fd_sc_hd__clkbuf_16 \Tile_X0Y1_DSP_bot/strobe_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[6] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/strobe_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[7] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/strobe_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[8] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Tile_X0Y1_FrameStrobe_O[9] ));
 sky130_fd_sc_hd__buf_4 input1 (.A(Tile_X0Y0_E1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(Tile_X0Y0_E2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(Tile_X0Y0_S2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(Tile_X0Y0_S4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(Tile_X0Y0_S4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(Tile_X0Y0_S4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(Tile_X0Y0_S4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(Tile_X0Y0_S4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(Tile_X0Y0_S4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(Tile_X0Y0_S4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(Tile_X0Y0_S4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(Tile_X0Y0_S4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input11 (.A(Tile_X0Y0_E2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(Tile_X0Y0_S4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(Tile_X0Y0_S4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(Tile_X0Y0_S4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(Tile_X0Y0_S4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(Tile_X0Y0_S4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(Tile_X0Y0_S4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(Tile_X0Y0_S4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(Tile_X0Y0_SS4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(Tile_X0Y0_SS4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(Tile_X0Y0_SS4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input12 (.A(Tile_X0Y0_E2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(Tile_X0Y0_SS4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(Tile_X0Y0_SS4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(Tile_X0Y0_SS4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(Tile_X0Y0_SS4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__buf_2 input124 (.A(Tile_X0Y0_SS4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(Tile_X0Y0_SS4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input126 (.A(Tile_X0Y0_SS4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(Tile_X0Y0_SS4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__buf_1 input128 (.A(Tile_X0Y0_SS4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(Tile_X0Y0_SS4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input13 (.A(Tile_X0Y0_E2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(Tile_X0Y0_SS4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(Tile_X0Y0_SS4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(Tile_X0Y0_SS4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__buf_4 input133 (.A(Tile_X0Y0_W1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__buf_4 input134 (.A(Tile_X0Y0_W1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__buf_4 input135 (.A(Tile_X0Y0_W1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__buf_4 input136 (.A(Tile_X0Y0_W1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(Tile_X0Y0_W2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(Tile_X0Y0_W2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(Tile_X0Y0_W2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(Tile_X0Y0_E2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input140 (.A(Tile_X0Y0_W2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 input141 (.A(Tile_X0Y0_W2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(Tile_X0Y0_W2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 input143 (.A(Tile_X0Y0_W2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 input144 (.A(Tile_X0Y0_W2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input145 (.A(Tile_X0Y0_W2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__buf_2 input146 (.A(Tile_X0Y0_W2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__buf_2 input147 (.A(Tile_X0Y0_W2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 input148 (.A(Tile_X0Y0_W2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(Tile_X0Y0_W2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__buf_2 input15 (.A(Tile_X0Y0_E2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input150 (.A(Tile_X0Y0_W2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 input151 (.A(Tile_X0Y0_W2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 input152 (.A(Tile_X0Y0_W2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(Tile_X0Y0_W6END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(Tile_X0Y0_W6END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(Tile_X0Y0_W6END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__buf_4 input156 (.A(Tile_X0Y0_W6END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(Tile_X0Y0_W6END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(Tile_X0Y0_W6END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(Tile_X0Y0_W6END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__buf_2 input16 (.A(Tile_X0Y0_E2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(Tile_X0Y0_W6END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(Tile_X0Y0_W6END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(Tile_X0Y0_W6END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(Tile_X0Y0_W6END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(Tile_X0Y0_W6END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 input165 (.A(Tile_X0Y0_WW4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(Tile_X0Y0_WW4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(Tile_X0Y0_WW4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(Tile_X0Y0_WW4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(Tile_X0Y0_WW4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(Tile_X0Y0_E2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(Tile_X0Y0_WW4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(Tile_X0Y0_WW4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(Tile_X0Y0_WW4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(Tile_X0Y0_WW4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 input174 (.A(Tile_X0Y0_WW4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(Tile_X0Y0_WW4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(Tile_X0Y0_WW4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(Tile_X0Y0_WW4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(Tile_X0Y0_WW4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(Tile_X0Y0_WW4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(Tile_X0Y0_E2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(Tile_X0Y0_WW4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 input181 (.A(Tile_X0Y1_E1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 input182 (.A(Tile_X0Y1_E1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 input183 (.A(Tile_X0Y1_E1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__buf_4 input184 (.A(Tile_X0Y1_E1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__buf_2 input185 (.A(Tile_X0Y1_E2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(Tile_X0Y1_E2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 input187 (.A(Tile_X0Y1_E2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 input188 (.A(Tile_X0Y1_E2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 input189 (.A(Tile_X0Y1_E2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__buf_2 input19 (.A(Tile_X0Y0_E2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(Tile_X0Y1_E2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(Tile_X0Y1_E2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 input192 (.A(Tile_X0Y1_E2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__buf_2 input193 (.A(Tile_X0Y1_E2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__buf_2 input194 (.A(Tile_X0Y1_E2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__buf_2 input195 (.A(Tile_X0Y1_E2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__buf_2 input196 (.A(Tile_X0Y1_E2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__buf_2 input197 (.A(Tile_X0Y1_E2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 input198 (.A(Tile_X0Y1_E2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 input199 (.A(Tile_X0Y1_E2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__buf_4 input2 (.A(Tile_X0Y0_E1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(Tile_X0Y0_E2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input200 (.A(Tile_X0Y1_E2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__buf_4 input201 (.A(Tile_X0Y1_E6END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(Tile_X0Y1_E6END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(Tile_X0Y1_E6END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__buf_4 input204 (.A(Tile_X0Y1_E6END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(Tile_X0Y1_E6END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 input206 (.A(Tile_X0Y1_E6END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 input207 (.A(Tile_X0Y1_E6END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(Tile_X0Y1_E6END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(Tile_X0Y1_E6END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__buf_4 input21 (.A(Tile_X0Y0_E6END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(Tile_X0Y1_E6END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(Tile_X0Y1_E6END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(Tile_X0Y1_E6END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(Tile_X0Y1_EE4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(Tile_X0Y1_EE4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(Tile_X0Y1_EE4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(Tile_X0Y1_EE4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 input217 (.A(Tile_X0Y1_EE4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(Tile_X0Y1_EE4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 input219 (.A(Tile_X0Y1_EE4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(Tile_X0Y0_E6END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input220 (.A(Tile_X0Y1_EE4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 input221 (.A(Tile_X0Y1_EE4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__buf_1 input222 (.A(Tile_X0Y1_EE4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(Tile_X0Y1_EE4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 input224 (.A(Tile_X0Y1_EE4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 input225 (.A(Tile_X0Y1_EE4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 input226 (.A(Tile_X0Y1_EE4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(Tile_X0Y1_EE4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(Tile_X0Y1_EE4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 input229 (.A(Tile_X0Y1_FrameData[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(Tile_X0Y0_E6END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_8 input230 (.A(Tile_X0Y1_FrameData[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 input231 (.A(Tile_X0Y1_FrameData[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_8 input232 (.A(Tile_X0Y1_FrameData[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_8 input233 (.A(Tile_X0Y1_FrameData[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_8 input234 (.A(Tile_X0Y1_FrameData[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_8 input235 (.A(Tile_X0Y1_FrameData[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net235));
 sky130_fd_sc_hd__buf_4 input236 (.A(Tile_X0Y1_FrameData[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net236));
 sky130_fd_sc_hd__buf_4 input237 (.A(Tile_X0Y1_FrameData[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_8 input238 (.A(Tile_X0Y1_FrameData[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_8 input239 (.A(Tile_X0Y1_FrameData[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net239));
 sky130_fd_sc_hd__buf_4 input24 (.A(Tile_X0Y0_E6END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_8 input240 (.A(Tile_X0Y1_FrameData[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_8 input241 (.A(Tile_X0Y1_FrameData[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_8 input242 (.A(Tile_X0Y1_FrameData[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_8 input243 (.A(Tile_X0Y1_FrameData[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_8 input244 (.A(Tile_X0Y1_FrameData[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net244));
 sky130_fd_sc_hd__buf_4 input245 (.A(Tile_X0Y1_FrameData[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net245));
 sky130_fd_sc_hd__buf_4 input246 (.A(Tile_X0Y1_FrameData[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_8 input247 (.A(Tile_X0Y1_FrameData[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_8 input248 (.A(Tile_X0Y1_FrameData[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_8 input249 (.A(Tile_X0Y1_FrameData[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(Tile_X0Y0_E6END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__buf_6 input250 (.A(Tile_X0Y1_FrameData[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net250));
 sky130_fd_sc_hd__buf_6 input251 (.A(Tile_X0Y1_FrameData[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net251));
 sky130_fd_sc_hd__buf_6 input252 (.A(Tile_X0Y1_FrameData[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 input253 (.A(Tile_X0Y1_FrameData[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net253));
 sky130_fd_sc_hd__buf_6 input254 (.A(Tile_X0Y1_FrameData[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net254));
 sky130_fd_sc_hd__buf_6 input255 (.A(Tile_X0Y1_FrameData[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net255));
 sky130_fd_sc_hd__buf_6 input256 (.A(Tile_X0Y1_FrameData[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_8 input257 (.A(Tile_X0Y1_FrameData[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net257));
 sky130_fd_sc_hd__buf_6 input258 (.A(Tile_X0Y1_FrameData[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_8 input259 (.A(Tile_X0Y1_FrameData[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(Tile_X0Y0_E6END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_8 input260 (.A(Tile_X0Y1_FrameData[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net260));
 sky130_fd_sc_hd__buf_8 input261 (.A(Tile_X0Y1_FrameStrobe[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net261));
 sky130_fd_sc_hd__buf_8 input262 (.A(Tile_X0Y1_FrameStrobe[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net262));
 sky130_fd_sc_hd__buf_8 input263 (.A(Tile_X0Y1_FrameStrobe[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net263));
 sky130_fd_sc_hd__buf_12 input264 (.A(Tile_X0Y1_FrameStrobe[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 input265 (.A(Tile_X0Y1_FrameStrobe[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 input266 (.A(Tile_X0Y1_FrameStrobe[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 input267 (.A(Tile_X0Y1_FrameStrobe[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 input268 (.A(Tile_X0Y1_FrameStrobe[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 input269 (.A(Tile_X0Y1_FrameStrobe[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(Tile_X0Y0_E6END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input270 (.A(Tile_X0Y1_FrameStrobe[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 input271 (.A(Tile_X0Y1_FrameStrobe[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net271));
 sky130_fd_sc_hd__buf_12 input272 (.A(Tile_X0Y1_FrameStrobe[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net272));
 sky130_fd_sc_hd__buf_8 input273 (.A(Tile_X0Y1_FrameStrobe[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net273));
 sky130_fd_sc_hd__buf_12 input274 (.A(Tile_X0Y1_FrameStrobe[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_16 input275 (.A(Tile_X0Y1_FrameStrobe[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_16 input276 (.A(Tile_X0Y1_FrameStrobe[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_16 input277 (.A(Tile_X0Y1_FrameStrobe[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net277));
 sky130_fd_sc_hd__buf_8 input278 (.A(Tile_X0Y1_FrameStrobe[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net278));
 sky130_fd_sc_hd__buf_8 input279 (.A(Tile_X0Y1_FrameStrobe[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(Tile_X0Y0_E6END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_16 input280 (.A(Tile_X0Y1_FrameStrobe[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net280));
 sky130_fd_sc_hd__buf_4 input281 (.A(Tile_X0Y1_N1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net281));
 sky130_fd_sc_hd__buf_4 input282 (.A(Tile_X0Y1_N1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 input283 (.A(Tile_X0Y1_N1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_4 input284 (.A(Tile_X0Y1_N1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 input285 (.A(Tile_X0Y1_N2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 input286 (.A(Tile_X0Y1_N2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 input287 (.A(Tile_X0Y1_N2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net287));
 sky130_fd_sc_hd__buf_2 input288 (.A(Tile_X0Y1_N2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 input289 (.A(Tile_X0Y1_N2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(Tile_X0Y0_E6END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input290 (.A(Tile_X0Y1_N2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net290));
 sky130_fd_sc_hd__buf_2 input291 (.A(Tile_X0Y1_N2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net291));
 sky130_fd_sc_hd__buf_2 input292 (.A(Tile_X0Y1_N2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net292));
 sky130_fd_sc_hd__buf_2 input293 (.A(Tile_X0Y1_N2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net293));
 sky130_fd_sc_hd__buf_2 input294 (.A(Tile_X0Y1_N2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 input295 (.A(Tile_X0Y1_N2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 input296 (.A(Tile_X0Y1_N2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net296));
 sky130_fd_sc_hd__buf_2 input297 (.A(Tile_X0Y1_N2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net297));
 sky130_fd_sc_hd__buf_2 input298 (.A(Tile_X0Y1_N2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net298));
 sky130_fd_sc_hd__buf_4 input299 (.A(Tile_X0Y1_N2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net299));
 sky130_fd_sc_hd__buf_4 input3 (.A(Tile_X0Y0_E1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(Tile_X0Y0_E6END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input300 (.A(Tile_X0Y1_N2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 input301 (.A(Tile_X0Y1_N4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 input302 (.A(Tile_X0Y1_N4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 input303 (.A(Tile_X0Y1_N4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 input304 (.A(Tile_X0Y1_N4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 input305 (.A(Tile_X0Y1_N4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 input306 (.A(Tile_X0Y1_N4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 input307 (.A(Tile_X0Y1_N4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net307));
 sky130_fd_sc_hd__dlymetal6s2s_1 input308 (.A(Tile_X0Y1_N4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 input309 (.A(Tile_X0Y1_N4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(Tile_X0Y0_E6END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input310 (.A(Tile_X0Y1_N4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 input311 (.A(Tile_X0Y1_N4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 input312 (.A(Tile_X0Y1_N4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 input313 (.A(Tile_X0Y1_N4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 input314 (.A(Tile_X0Y1_N4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 input315 (.A(Tile_X0Y1_N4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 input316 (.A(Tile_X0Y1_N4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net316));
 sky130_fd_sc_hd__buf_1 input317 (.A(Tile_X0Y1_NN4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 input318 (.A(Tile_X0Y1_NN4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 input319 (.A(Tile_X0Y1_NN4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(Tile_X0Y0_E6END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input320 (.A(Tile_X0Y1_NN4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 input321 (.A(Tile_X0Y1_NN4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 input322 (.A(Tile_X0Y1_NN4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 input323 (.A(Tile_X0Y1_NN4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 input324 (.A(Tile_X0Y1_NN4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 input325 (.A(Tile_X0Y1_NN4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 input326 (.A(Tile_X0Y1_NN4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 input327 (.A(Tile_X0Y1_NN4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 input328 (.A(Tile_X0Y1_NN4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 input329 (.A(Tile_X0Y1_NN4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net329));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(Tile_X0Y0_EE4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input330 (.A(Tile_X0Y1_NN4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 input331 (.A(Tile_X0Y1_NN4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 input332 (.A(Tile_X0Y1_NN4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net332));
 sky130_fd_sc_hd__buf_12 input333 (.A(Tile_X0Y1_UserCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 input334 (.A(Tile_X0Y1_W1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net334));
 sky130_fd_sc_hd__buf_4 input335 (.A(Tile_X0Y1_W1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net335));
 sky130_fd_sc_hd__buf_4 input336 (.A(Tile_X0Y1_W1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net336));
 sky130_fd_sc_hd__buf_4 input337 (.A(Tile_X0Y1_W1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net337));
 sky130_fd_sc_hd__buf_2 input338 (.A(Tile_X0Y1_W2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net338));
 sky130_fd_sc_hd__buf_2 input339 (.A(Tile_X0Y1_W2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(Tile_X0Y0_EE4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input340 (.A(Tile_X0Y1_W2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 input341 (.A(Tile_X0Y1_W2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 input342 (.A(Tile_X0Y1_W2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 input343 (.A(Tile_X0Y1_W2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net343));
 sky130_fd_sc_hd__dlymetal6s2s_1 input344 (.A(Tile_X0Y1_W2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 input345 (.A(Tile_X0Y1_W2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 input346 (.A(Tile_X0Y1_W2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net346));
 sky130_fd_sc_hd__buf_2 input347 (.A(Tile_X0Y1_W2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_4 input348 (.A(Tile_X0Y1_W2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_4 input349 (.A(Tile_X0Y1_W2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(Tile_X0Y0_EE4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input350 (.A(Tile_X0Y1_W2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_4 input351 (.A(Tile_X0Y1_W2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_4 input352 (.A(Tile_X0Y1_W2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_4 input353 (.A(Tile_X0Y1_W2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 input354 (.A(Tile_X0Y1_W6END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 input355 (.A(Tile_X0Y1_W6END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 input356 (.A(Tile_X0Y1_W6END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_4 input357 (.A(Tile_X0Y1_W6END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 input358 (.A(Tile_X0Y1_W6END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 input359 (.A(Tile_X0Y1_W6END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(Tile_X0Y0_EE4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input360 (.A(Tile_X0Y1_W6END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 input361 (.A(Tile_X0Y1_W6END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 input362 (.A(Tile_X0Y1_W6END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 input363 (.A(Tile_X0Y1_W6END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 input364 (.A(Tile_X0Y1_W6END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 input365 (.A(Tile_X0Y1_W6END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net365));
 sky130_fd_sc_hd__buf_2 input366 (.A(Tile_X0Y1_WW4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 input367 (.A(Tile_X0Y1_WW4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 input368 (.A(Tile_X0Y1_WW4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 input369 (.A(Tile_X0Y1_WW4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(Tile_X0Y0_EE4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input370 (.A(Tile_X0Y1_WW4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 input371 (.A(Tile_X0Y1_WW4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 input372 (.A(Tile_X0Y1_WW4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 input373 (.A(Tile_X0Y1_WW4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net373));
 sky130_fd_sc_hd__buf_2 input374 (.A(Tile_X0Y1_WW4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net374));
 sky130_fd_sc_hd__dlymetal6s2s_1 input375 (.A(Tile_X0Y1_WW4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 input376 (.A(Tile_X0Y1_WW4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 input377 (.A(Tile_X0Y1_WW4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 input378 (.A(Tile_X0Y1_WW4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 input379 (.A(Tile_X0Y1_WW4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(Tile_X0Y0_EE4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input380 (.A(Tile_X0Y1_WW4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 input381 (.A(Tile_X0Y1_WW4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(Tile_X0Y0_EE4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(Tile_X0Y0_E1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(Tile_X0Y0_EE4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(Tile_X0Y0_EE4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(Tile_X0Y0_EE4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(Tile_X0Y0_EE4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(Tile_X0Y0_EE4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(Tile_X0Y0_EE4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(Tile_X0Y0_EE4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(Tile_X0Y0_EE4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(Tile_X0Y0_EE4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 input49 (.A(Tile_X0Y0_FrameData[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(Tile_X0Y0_E2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input50 (.A(Tile_X0Y0_FrameData[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 input51 (.A(Tile_X0Y0_FrameData[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_8 input52 (.A(Tile_X0Y0_FrameData[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_8 input53 (.A(Tile_X0Y0_FrameData[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_6 input54 (.A(Tile_X0Y0_FrameData[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 input55 (.A(Tile_X0Y0_FrameData[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 input56 (.A(Tile_X0Y0_FrameData[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(Tile_X0Y0_FrameData[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__buf_6 input58 (.A(Tile_X0Y0_FrameData[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__buf_6 input59 (.A(Tile_X0Y0_FrameData[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input6 (.A(Tile_X0Y0_E2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 input60 (.A(Tile_X0Y0_FrameData[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(Tile_X0Y0_FrameData[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 input62 (.A(Tile_X0Y0_FrameData[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__buf_6 input63 (.A(Tile_X0Y0_FrameData[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 input64 (.A(Tile_X0Y0_FrameData[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_8 input65 (.A(Tile_X0Y0_FrameData[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_8 input66 (.A(Tile_X0Y0_FrameData[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input67 (.A(Tile_X0Y0_FrameData[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_8 input68 (.A(Tile_X0Y0_FrameData[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__buf_6 input69 (.A(Tile_X0Y0_FrameData[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input7 (.A(Tile_X0Y0_E2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input70 (.A(Tile_X0Y0_FrameData[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_8 input71 (.A(Tile_X0Y0_FrameData[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 input72 (.A(Tile_X0Y0_FrameData[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_8 input73 (.A(Tile_X0Y0_FrameData[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_8 input74 (.A(Tile_X0Y0_FrameData[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__buf_6 input75 (.A(Tile_X0Y0_FrameData[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__buf_6 input76 (.A(Tile_X0Y0_FrameData[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_8 input77 (.A(Tile_X0Y0_FrameData[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_8 input78 (.A(Tile_X0Y0_FrameData[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(Tile_X0Y0_FrameData[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(Tile_X0Y0_E2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input80 (.A(Tile_X0Y0_FrameData[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(Tile_X0Y0_S1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(Tile_X0Y0_S1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(Tile_X0Y0_S1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(Tile_X0Y0_S1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input85 (.A(Tile_X0Y0_S2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 input86 (.A(Tile_X0Y0_S2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(Tile_X0Y0_S2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(Tile_X0Y0_S2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(Tile_X0Y0_S2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(Tile_X0Y0_E2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input90 (.A(Tile_X0Y0_S2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(Tile_X0Y0_S2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(Tile_X0Y0_S2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(Tile_X0Y0_S2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(Tile_X0Y0_S2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 input95 (.A(Tile_X0Y0_S2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__buf_4 input96 (.A(Tile_X0Y0_S2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__buf_4 input97 (.A(Tile_X0Y0_S2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(Tile_X0Y0_S2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 input99 (.A(Tile_X0Y0_S2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__buf_12 max_cap763 (.A(\Tile_X0Y1_DSP_bot/Q6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_8 max_cap764 (.A(\Tile_X0Y1_DSP_bot/Q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net764));
 sky130_fd_sc_hd__buf_2 output382 (.A(net382),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E1BEG[0]));
 sky130_fd_sc_hd__buf_2 output383 (.A(net383),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output385 (.A(net385),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E1BEG[3]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEG[0]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net387),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output389 (.A(net389),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output390 (.A(net390),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output391 (.A(net391),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEG[5]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEG[6]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net393),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output394 (.A(net394),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output395 (.A(net395),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output397 (.A(net397),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output398 (.A(net398),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output399 (.A(net399),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output400 (.A(net400),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output401 (.A(net401),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output402 (.A(net402),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output403 (.A(net403),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output404 (.A(net404),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net405),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output406 (.A(net406),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output407 (.A(net407),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output408 (.A(net408),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net409),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output410 (.A(net410),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output411 (.A(net411),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output412 (.A(net412),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output413 (.A(net413),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output414 (.A(net414),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output416 (.A(net416),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output417 (.A(net417),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output418 (.A(net418),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net419),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[14]));
 sky130_fd_sc_hd__buf_2 output420 (.A(net420),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output421 (.A(net421),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output422 (.A(net422),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output423 (.A(net423),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output424 (.A(net424),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output425 (.A(net425),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output426 (.A(net426),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output427 (.A(net427),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output428 (.A(net428),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output429 (.A(net429),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_EE4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output430 (.A(net430),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output431 (.A(net431),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output432 (.A(net432),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net433),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output434 (.A(net434),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output435 (.A(net435),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output436 (.A(net436),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output437 (.A(net437),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output438 (.A(net438),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output439 (.A(net439),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output440 (.A(net440),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output441 (.A(net441),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output442 (.A(net442),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output443 (.A(net443),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output444 (.A(net444),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output445 (.A(net445),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output446 (.A(net446),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[24]));
 sky130_fd_sc_hd__clkbuf_4 output447 (.A(net447),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[25]));
 sky130_fd_sc_hd__clkbuf_4 output448 (.A(net448),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output449 (.A(net449),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output450 (.A(net450),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output451 (.A(net451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output452 (.A(net452),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output453 (.A(net453),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output454 (.A(net454),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output455 (.A(net455),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output456 (.A(net456),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output457 (.A(net457),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output458 (.A(net458),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output459 (.A(net459),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output460 (.A(net460),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output461 (.A(net461),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameData_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output462 (.A(net462),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output463 (.A(net463),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output464 (.A(net464),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output465 (.A(net465),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output466 (.A(net466),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output467 (.A(net467),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output468 (.A(net468),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output469 (.A(net469),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output470 (.A(net470),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output471 (.A(net471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output472 (.A(net472),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output473 (.A(net473),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output474 (.A(net474),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output475 (.A(net475),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output476 (.A(net476),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output477 (.A(net477),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output478 (.A(net478),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output479 (.A(net479),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output480 (.A(net480),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output481 (.A(net481),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_FrameStrobe_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output482 (.A(net482),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output483 (.A(net483),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output484 (.A(net484),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output485 (.A(net485),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output486 (.A(net486),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output487 (.A(net487),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output488 (.A(net488),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output489 (.A(net489),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output490 (.A(net490),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output491 (.A(net491),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output492 (.A(net492),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output493 (.A(net493),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output494 (.A(net494),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output495 (.A(net495),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output496 (.A(net496),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output497 (.A(net497),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output498 (.A(net498),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output499 (.A(net499),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output500 (.A(net500),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output501 (.A(net501),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output502 (.A(net502),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output503 (.A(net503),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output504 (.A(net504),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output505 (.A(net505),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output506 (.A(net506),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output507 (.A(net507),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output508 (.A(net508),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output509 (.A(net509),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output510 (.A(net510),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output511 (.A(net511),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output512 (.A(net512),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output513 (.A(net513),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output514 (.A(net514),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output515 (.A(net515),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output516 (.A(net516),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output517 (.A(net517),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_N4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output518 (.A(net518),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output519 (.A(net519),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output520 (.A(net520),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output521 (.A(net521),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output522 (.A(net522),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output523 (.A(net523),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output524 (.A(net524),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output525 (.A(net525),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output526 (.A(net526),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output527 (.A(net527),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output528 (.A(net528),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output529 (.A(net529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output530 (.A(net530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output531 (.A(net531),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output532 (.A(net532),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output533 (.A(net533),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_NN4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output534 (.A(net534),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output535 (.A(net535),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output536 (.A(net536),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output537 (.A(net537),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output538 (.A(net538),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output539 (.A(net539),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output540 (.A(net540),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output541 (.A(net541),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output542 (.A(net542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output543 (.A(net543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output544 (.A(net544),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output545 (.A(net545),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output546 (.A(net546),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output547 (.A(net547),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output548 (.A(net548),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output549 (.A(net549),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output550 (.A(net550),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output551 (.A(net551),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output552 (.A(net552),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output553 (.A(net553),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output554 (.A(net554),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output555 (.A(net555),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output556 (.A(net556),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output557 (.A(net557),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output558 (.A(net558),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output559 (.A(net559),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output560 (.A(net560),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output561 (.A(net561),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output562 (.A(net562),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output563 (.A(net563),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output564 (.A(net564),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output565 (.A(net565),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output566 (.A(net566),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_W6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output567 (.A(net567),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output568 (.A(net568),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output569 (.A(net569),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output570 (.A(net570),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output571 (.A(net571),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output572 (.A(net572),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output573 (.A(net573),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output574 (.A(net574),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output575 (.A(net575),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output576 (.A(net576),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output577 (.A(net577),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output578 (.A(net578),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output579 (.A(net579),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output580 (.A(net580),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output581 (.A(net581),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output582 (.A(net582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y0_WW4BEG[9]));
 sky130_fd_sc_hd__buf_2 output583 (.A(net583),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E1BEG[0]));
 sky130_fd_sc_hd__buf_2 output584 (.A(net584),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output585 (.A(net585),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output586 (.A(net586),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output587 (.A(net587),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output588 (.A(net588),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output589 (.A(net589),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output590 (.A(net590),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output591 (.A(net591),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output592 (.A(net592),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output593 (.A(net593),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output594 (.A(net594),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output595 (.A(net595),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output596 (.A(net596),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output597 (.A(net597),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output598 (.A(net598),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output599 (.A(net599),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output600 (.A(net600),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output601 (.A(net601),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output602 (.A(net602),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output603 (.A(net603),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output604 (.A(net604),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output605 (.A(net605),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output606 (.A(net606),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output607 (.A(net607),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output608 (.A(net608),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output609 (.A(net609),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output610 (.A(net610),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output611 (.A(net611),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output612 (.A(net612),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output613 (.A(net613),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output614 (.A(net614),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_E6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output615 (.A(net615),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output616 (.A(net616),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output617 (.A(net617),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output618 (.A(net618),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[12]));
 sky130_fd_sc_hd__buf_2 output619 (.A(net619),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output620 (.A(net620),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output621 (.A(net621),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output622 (.A(net622),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output623 (.A(net623),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output624 (.A(net624),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output625 (.A(net625),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output626 (.A(net626),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output627 (.A(net627),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output628 (.A(net628),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output629 (.A(net629),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output630 (.A(net630),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output631 (.A(net631),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output632 (.A(net632),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output633 (.A(net633),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output634 (.A(net634),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output635 (.A(net635),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output636 (.A(net636),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output637 (.A(net637),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output638 (.A(net638),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output639 (.A(net639),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output640 (.A(net640),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output641 (.A(net641),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output642 (.A(net642),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output643 (.A(net643),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output644 (.A(net644),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output645 (.A(net645),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[22]));
 sky130_fd_sc_hd__clkbuf_4 output646 (.A(net646),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output647 (.A(net647),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output648 (.A(net648),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output649 (.A(net649),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output650 (.A(net650),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[27]));
 sky130_fd_sc_hd__clkbuf_4 output651 (.A(net651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output652 (.A(net652),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[29]));
 sky130_fd_sc_hd__clkbuf_4 output653 (.A(net653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output654 (.A(net654),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output655 (.A(net655),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[31]));
 sky130_fd_sc_hd__clkbuf_4 output656 (.A(net656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output657 (.A(net657),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output658 (.A(net658),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output659 (.A(net659),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output660 (.A(net660),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output661 (.A(net661),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output662 (.A(net662),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output663 (.A(net663),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output664 (.A(net664),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output665 (.A(net665),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output666 (.A(net666),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output667 (.A(net667),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output668 (.A(net668),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output669 (.A(net669),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output670 (.A(net670),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output671 (.A(net671),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output672 (.A(net672),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output673 (.A(net673),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output674 (.A(net674),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output675 (.A(net675),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output676 (.A(net676),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output677 (.A(net677),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output678 (.A(net678),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output679 (.A(net679),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output680 (.A(net680),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output681 (.A(net681),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output682 (.A(net682),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output683 (.A(net683),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output684 (.A(net684),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output685 (.A(net685),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output686 (.A(net686),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output687 (.A(net687),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output688 (.A(net688),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output689 (.A(net689),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output690 (.A(net690),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output691 (.A(net691),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output692 (.A(net692),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output693 (.A(net693),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output694 (.A(net694),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output695 (.A(net695),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output696 (.A(net696),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output697 (.A(net697),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output698 (.A(net698),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output699 (.A(net699),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output700 (.A(net700),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output701 (.A(net701),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output702 (.A(net702),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output703 (.A(net703),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output704 (.A(net704),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output705 (.A(net705),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output706 (.A(net706),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output707 (.A(net707),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output708 (.A(net708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output709 (.A(net709),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output710 (.A(net710),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output711 (.A(net711),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output712 (.A(net712),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output713 (.A(net713),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[8]));
 sky130_fd_sc_hd__buf_2 output714 (.A(net714),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_SS4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output715 (.A(net715),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output716 (.A(net716),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output717 (.A(net717),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output718 (.A(net718),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output719 (.A(net719),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output720 (.A(net720),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output721 (.A(net721),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output722 (.A(net722),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output723 (.A(net723),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output724 (.A(net724),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output725 (.A(net725),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output726 (.A(net726),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output727 (.A(net727),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output728 (.A(net728),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output729 (.A(net729),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output730 (.A(net730),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output731 (.A(net731),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output732 (.A(net732),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output733 (.A(net733),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output734 (.A(net734),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output735 (.A(net735),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output736 (.A(net736),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output737 (.A(net737),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output738 (.A(net738),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output739 (.A(net739),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output740 (.A(net740),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output741 (.A(net741),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output742 (.A(net742),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output743 (.A(net743),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output744 (.A(net744),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output745 (.A(net745),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output746 (.A(net746),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_W6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output747 (.A(net747),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output748 (.A(net748),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output749 (.A(net749),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output750 (.A(net750),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output751 (.A(net751),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output752 (.A(net752),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output753 (.A(net753),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output754 (.A(net754),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output755 (.A(net755),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output756 (.A(net756),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output757 (.A(net757),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output758 (.A(net758),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output759 (.A(net759),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output760 (.A(net760),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output761 (.A(net761),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output762 (.A(net762),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Tile_X0Y1_WW4BEG[9]));
endmodule
