magic
tech sky130A
magscale 1 2
timestamp 1733394402
<< obsli1 >>
rect 1104 1071 45816 8721
<< obsm1 >>
rect 658 620 46354 9988
<< metal2 >>
rect 662 9840 718 10000
rect 1030 9840 1086 10000
rect 1398 9840 1454 10000
rect 1766 9840 1822 10000
rect 2134 9840 2190 10000
rect 2502 9840 2558 10000
rect 2870 9840 2926 10000
rect 3238 9840 3294 10000
rect 3606 9840 3662 10000
rect 3974 9840 4030 10000
rect 4342 9840 4398 10000
rect 4710 9840 4766 10000
rect 5078 9840 5134 10000
rect 5446 9840 5502 10000
rect 5814 9840 5870 10000
rect 6182 9840 6238 10000
rect 6550 9840 6606 10000
rect 6918 9840 6974 10000
rect 7286 9840 7342 10000
rect 7654 9840 7710 10000
rect 8022 9840 8078 10000
rect 8390 9840 8446 10000
rect 8758 9840 8814 10000
rect 9126 9840 9182 10000
rect 9494 9840 9550 10000
rect 9862 9840 9918 10000
rect 10230 9840 10286 10000
rect 10598 9840 10654 10000
rect 10966 9840 11022 10000
rect 11334 9840 11390 10000
rect 11702 9840 11758 10000
rect 12070 9840 12126 10000
rect 12438 9840 12494 10000
rect 12806 9840 12862 10000
rect 13174 9840 13230 10000
rect 13542 9840 13598 10000
rect 13910 9840 13966 10000
rect 14278 9840 14334 10000
rect 14646 9840 14702 10000
rect 15014 9840 15070 10000
rect 15382 9840 15438 10000
rect 15750 9840 15806 10000
rect 16118 9840 16174 10000
rect 16486 9840 16542 10000
rect 16854 9840 16910 10000
rect 17222 9840 17278 10000
rect 17590 9840 17646 10000
rect 17958 9840 18014 10000
rect 18326 9840 18382 10000
rect 18694 9840 18750 10000
rect 19062 9840 19118 10000
rect 19430 9840 19486 10000
rect 19798 9840 19854 10000
rect 20166 9840 20222 10000
rect 20534 9840 20590 10000
rect 20902 9840 20958 10000
rect 21270 9840 21326 10000
rect 21638 9840 21694 10000
rect 22006 9840 22062 10000
rect 22374 9840 22430 10000
rect 22742 9840 22798 10000
rect 23110 9840 23166 10000
rect 23478 9840 23534 10000
rect 23846 9840 23902 10000
rect 24214 9840 24270 10000
rect 24582 9840 24638 10000
rect 24950 9840 25006 10000
rect 25318 9840 25374 10000
rect 25686 9840 25742 10000
rect 26054 9840 26110 10000
rect 26422 9840 26478 10000
rect 26790 9840 26846 10000
rect 27158 9840 27214 10000
rect 27526 9840 27582 10000
rect 27894 9840 27950 10000
rect 28262 9840 28318 10000
rect 28630 9840 28686 10000
rect 28998 9840 29054 10000
rect 29366 9840 29422 10000
rect 29734 9840 29790 10000
rect 30102 9840 30158 10000
rect 30470 9840 30526 10000
rect 30838 9840 30894 10000
rect 31206 9840 31262 10000
rect 31574 9840 31630 10000
rect 31942 9840 31998 10000
rect 32310 9840 32366 10000
rect 32678 9840 32734 10000
rect 33046 9840 33102 10000
rect 33414 9840 33470 10000
rect 33782 9840 33838 10000
rect 34150 9840 34206 10000
rect 34518 9840 34574 10000
rect 34886 9840 34942 10000
rect 35254 9840 35310 10000
rect 35622 9840 35678 10000
rect 35990 9840 36046 10000
rect 36358 9840 36414 10000
rect 36726 9840 36782 10000
rect 37094 9840 37150 10000
rect 37462 9840 37518 10000
rect 37830 9840 37886 10000
rect 38198 9840 38254 10000
rect 38566 9840 38622 10000
rect 38934 9840 38990 10000
rect 39302 9840 39358 10000
rect 39670 9840 39726 10000
rect 40038 9840 40094 10000
rect 40406 9840 40462 10000
rect 40774 9840 40830 10000
rect 41142 9840 41198 10000
rect 41510 9840 41566 10000
rect 41878 9840 41934 10000
rect 42246 9840 42302 10000
rect 42614 9840 42670 10000
rect 42982 9840 43038 10000
rect 43350 9840 43406 10000
rect 43718 9840 43774 10000
rect 44086 9840 44142 10000
rect 44454 9840 44510 10000
rect 44822 9840 44878 10000
rect 45190 9840 45246 10000
rect 45558 9840 45614 10000
rect 45926 9840 45982 10000
rect 46294 9840 46350 10000
rect 1398 0 1454 160
rect 3606 0 3662 160
rect 5814 0 5870 160
rect 8022 0 8078 160
rect 10230 0 10286 160
rect 12438 0 12494 160
rect 14646 0 14702 160
rect 16854 0 16910 160
rect 19062 0 19118 160
rect 21270 0 21326 160
rect 23478 0 23534 160
rect 25686 0 25742 160
rect 27894 0 27950 160
rect 30102 0 30158 160
rect 32310 0 32366 160
rect 34518 0 34574 160
rect 36726 0 36782 160
rect 38934 0 38990 160
rect 41142 0 41198 160
rect 43350 0 43406 160
rect 45558 0 45614 160
<< obsm2 >>
rect 774 9784 974 9994
rect 1142 9784 1342 9994
rect 1510 9784 1710 9994
rect 1878 9784 2078 9994
rect 2246 9784 2446 9994
rect 2614 9784 2814 9994
rect 2982 9784 3182 9994
rect 3350 9784 3550 9994
rect 3718 9784 3918 9994
rect 4086 9784 4286 9994
rect 4454 9784 4654 9994
rect 4822 9784 5022 9994
rect 5190 9784 5390 9994
rect 5558 9784 5758 9994
rect 5926 9784 6126 9994
rect 6294 9784 6494 9994
rect 6662 9784 6862 9994
rect 7030 9784 7230 9994
rect 7398 9784 7598 9994
rect 7766 9784 7966 9994
rect 8134 9784 8334 9994
rect 8502 9784 8702 9994
rect 8870 9784 9070 9994
rect 9238 9784 9438 9994
rect 9606 9784 9806 9994
rect 9974 9784 10174 9994
rect 10342 9784 10542 9994
rect 10710 9784 10910 9994
rect 11078 9784 11278 9994
rect 11446 9784 11646 9994
rect 11814 9784 12014 9994
rect 12182 9784 12382 9994
rect 12550 9784 12750 9994
rect 12918 9784 13118 9994
rect 13286 9784 13486 9994
rect 13654 9784 13854 9994
rect 14022 9784 14222 9994
rect 14390 9784 14590 9994
rect 14758 9784 14958 9994
rect 15126 9784 15326 9994
rect 15494 9784 15694 9994
rect 15862 9784 16062 9994
rect 16230 9784 16430 9994
rect 16598 9784 16798 9994
rect 16966 9784 17166 9994
rect 17334 9784 17534 9994
rect 17702 9784 17902 9994
rect 18070 9784 18270 9994
rect 18438 9784 18638 9994
rect 18806 9784 19006 9994
rect 19174 9784 19374 9994
rect 19542 9784 19742 9994
rect 19910 9784 20110 9994
rect 20278 9784 20478 9994
rect 20646 9784 20846 9994
rect 21014 9784 21214 9994
rect 21382 9784 21582 9994
rect 21750 9784 21950 9994
rect 22118 9784 22318 9994
rect 22486 9784 22686 9994
rect 22854 9784 23054 9994
rect 23222 9784 23422 9994
rect 23590 9784 23790 9994
rect 23958 9784 24158 9994
rect 24326 9784 24526 9994
rect 24694 9784 24894 9994
rect 25062 9784 25262 9994
rect 25430 9784 25630 9994
rect 25798 9784 25998 9994
rect 26166 9784 26366 9994
rect 26534 9784 26734 9994
rect 26902 9784 27102 9994
rect 27270 9784 27470 9994
rect 27638 9784 27838 9994
rect 28006 9784 28206 9994
rect 28374 9784 28574 9994
rect 28742 9784 28942 9994
rect 29110 9784 29310 9994
rect 29478 9784 29678 9994
rect 29846 9784 30046 9994
rect 30214 9784 30414 9994
rect 30582 9784 30782 9994
rect 30950 9784 31150 9994
rect 31318 9784 31518 9994
rect 31686 9784 31886 9994
rect 32054 9784 32254 9994
rect 32422 9784 32622 9994
rect 32790 9784 32990 9994
rect 33158 9784 33358 9994
rect 33526 9784 33726 9994
rect 33894 9784 34094 9994
rect 34262 9784 34462 9994
rect 34630 9784 34830 9994
rect 34998 9784 35198 9994
rect 35366 9784 35566 9994
rect 35734 9784 35934 9994
rect 36102 9784 36302 9994
rect 36470 9784 36670 9994
rect 36838 9784 37038 9994
rect 37206 9784 37406 9994
rect 37574 9784 37774 9994
rect 37942 9784 38142 9994
rect 38310 9784 38510 9994
rect 38678 9784 38878 9994
rect 39046 9784 39246 9994
rect 39414 9784 39614 9994
rect 39782 9784 39982 9994
rect 40150 9784 40350 9994
rect 40518 9784 40718 9994
rect 40886 9784 41086 9994
rect 41254 9784 41454 9994
rect 41622 9784 41822 9994
rect 41990 9784 42190 9994
rect 42358 9784 42558 9994
rect 42726 9784 42926 9994
rect 43094 9784 43294 9994
rect 43462 9784 43662 9994
rect 43830 9784 44030 9994
rect 44198 9784 44398 9994
rect 44566 9784 44766 9994
rect 44934 9784 45134 9994
rect 45302 9784 45502 9994
rect 45670 9784 45870 9994
rect 46038 9784 46238 9994
rect 664 216 46348 9784
rect 664 54 1342 216
rect 1510 54 3550 216
rect 3718 54 5758 216
rect 5926 54 7966 216
rect 8134 54 10174 216
rect 10342 54 12382 216
rect 12550 54 14590 216
rect 14758 54 16798 216
rect 16966 54 19006 216
rect 19174 54 21214 216
rect 21382 54 23422 216
rect 23590 54 25630 216
rect 25798 54 27838 216
rect 28006 54 30046 216
rect 30214 54 32254 216
rect 32422 54 34462 216
rect 34630 54 36670 216
rect 36838 54 38878 216
rect 39046 54 41086 216
rect 41254 54 43294 216
rect 43462 54 45502 216
rect 45670 54 46348 216
<< obsm3 >>
rect 2681 1055 45974 9893
<< metal4 >>
rect 6533 1040 6853 8752
rect 12122 1040 12442 8752
rect 17711 1040 18031 8752
rect 23300 1040 23620 8752
rect 28889 1040 29209 8752
rect 34478 1040 34798 8752
rect 40067 1040 40387 8752
rect 45656 1040 45976 8752
<< obsm4 >>
rect 20667 7787 20733 9213
<< labels >>
rlabel metal2 s 3606 0 3662 160 6 FrameStrobe[0]
port 1 nsew signal input
rlabel metal2 s 25686 0 25742 160 6 FrameStrobe[10]
port 2 nsew signal input
rlabel metal2 s 27894 0 27950 160 6 FrameStrobe[11]
port 3 nsew signal input
rlabel metal2 s 30102 0 30158 160 6 FrameStrobe[12]
port 4 nsew signal input
rlabel metal2 s 32310 0 32366 160 6 FrameStrobe[13]
port 5 nsew signal input
rlabel metal2 s 34518 0 34574 160 6 FrameStrobe[14]
port 6 nsew signal input
rlabel metal2 s 36726 0 36782 160 6 FrameStrobe[15]
port 7 nsew signal input
rlabel metal2 s 38934 0 38990 160 6 FrameStrobe[16]
port 8 nsew signal input
rlabel metal2 s 41142 0 41198 160 6 FrameStrobe[17]
port 9 nsew signal input
rlabel metal2 s 43350 0 43406 160 6 FrameStrobe[18]
port 10 nsew signal input
rlabel metal2 s 45558 0 45614 160 6 FrameStrobe[19]
port 11 nsew signal input
rlabel metal2 s 5814 0 5870 160 6 FrameStrobe[1]
port 12 nsew signal input
rlabel metal2 s 8022 0 8078 160 6 FrameStrobe[2]
port 13 nsew signal input
rlabel metal2 s 10230 0 10286 160 6 FrameStrobe[3]
port 14 nsew signal input
rlabel metal2 s 12438 0 12494 160 6 FrameStrobe[4]
port 15 nsew signal input
rlabel metal2 s 14646 0 14702 160 6 FrameStrobe[5]
port 16 nsew signal input
rlabel metal2 s 16854 0 16910 160 6 FrameStrobe[6]
port 17 nsew signal input
rlabel metal2 s 19062 0 19118 160 6 FrameStrobe[7]
port 18 nsew signal input
rlabel metal2 s 21270 0 21326 160 6 FrameStrobe[8]
port 19 nsew signal input
rlabel metal2 s 23478 0 23534 160 6 FrameStrobe[9]
port 20 nsew signal input
rlabel metal2 s 39302 9840 39358 10000 6 FrameStrobe_O[0]
port 21 nsew signal output
rlabel metal2 s 42982 9840 43038 10000 6 FrameStrobe_O[10]
port 22 nsew signal output
rlabel metal2 s 43350 9840 43406 10000 6 FrameStrobe_O[11]
port 23 nsew signal output
rlabel metal2 s 43718 9840 43774 10000 6 FrameStrobe_O[12]
port 24 nsew signal output
rlabel metal2 s 44086 9840 44142 10000 6 FrameStrobe_O[13]
port 25 nsew signal output
rlabel metal2 s 44454 9840 44510 10000 6 FrameStrobe_O[14]
port 26 nsew signal output
rlabel metal2 s 44822 9840 44878 10000 6 FrameStrobe_O[15]
port 27 nsew signal output
rlabel metal2 s 45190 9840 45246 10000 6 FrameStrobe_O[16]
port 28 nsew signal output
rlabel metal2 s 45558 9840 45614 10000 6 FrameStrobe_O[17]
port 29 nsew signal output
rlabel metal2 s 45926 9840 45982 10000 6 FrameStrobe_O[18]
port 30 nsew signal output
rlabel metal2 s 46294 9840 46350 10000 6 FrameStrobe_O[19]
port 31 nsew signal output
rlabel metal2 s 39670 9840 39726 10000 6 FrameStrobe_O[1]
port 32 nsew signal output
rlabel metal2 s 40038 9840 40094 10000 6 FrameStrobe_O[2]
port 33 nsew signal output
rlabel metal2 s 40406 9840 40462 10000 6 FrameStrobe_O[3]
port 34 nsew signal output
rlabel metal2 s 40774 9840 40830 10000 6 FrameStrobe_O[4]
port 35 nsew signal output
rlabel metal2 s 41142 9840 41198 10000 6 FrameStrobe_O[5]
port 36 nsew signal output
rlabel metal2 s 41510 9840 41566 10000 6 FrameStrobe_O[6]
port 37 nsew signal output
rlabel metal2 s 41878 9840 41934 10000 6 FrameStrobe_O[7]
port 38 nsew signal output
rlabel metal2 s 42246 9840 42302 10000 6 FrameStrobe_O[8]
port 39 nsew signal output
rlabel metal2 s 42614 9840 42670 10000 6 FrameStrobe_O[9]
port 40 nsew signal output
rlabel metal2 s 662 9840 718 10000 6 N1BEG[0]
port 41 nsew signal output
rlabel metal2 s 1030 9840 1086 10000 6 N1BEG[1]
port 42 nsew signal output
rlabel metal2 s 1398 9840 1454 10000 6 N1BEG[2]
port 43 nsew signal output
rlabel metal2 s 1766 9840 1822 10000 6 N1BEG[3]
port 44 nsew signal output
rlabel metal2 s 2134 9840 2190 10000 6 N2BEG[0]
port 45 nsew signal output
rlabel metal2 s 2502 9840 2558 10000 6 N2BEG[1]
port 46 nsew signal output
rlabel metal2 s 2870 9840 2926 10000 6 N2BEG[2]
port 47 nsew signal output
rlabel metal2 s 3238 9840 3294 10000 6 N2BEG[3]
port 48 nsew signal output
rlabel metal2 s 3606 9840 3662 10000 6 N2BEG[4]
port 49 nsew signal output
rlabel metal2 s 3974 9840 4030 10000 6 N2BEG[5]
port 50 nsew signal output
rlabel metal2 s 4342 9840 4398 10000 6 N2BEG[6]
port 51 nsew signal output
rlabel metal2 s 4710 9840 4766 10000 6 N2BEG[7]
port 52 nsew signal output
rlabel metal2 s 5078 9840 5134 10000 6 N2BEGb[0]
port 53 nsew signal output
rlabel metal2 s 5446 9840 5502 10000 6 N2BEGb[1]
port 54 nsew signal output
rlabel metal2 s 5814 9840 5870 10000 6 N2BEGb[2]
port 55 nsew signal output
rlabel metal2 s 6182 9840 6238 10000 6 N2BEGb[3]
port 56 nsew signal output
rlabel metal2 s 6550 9840 6606 10000 6 N2BEGb[4]
port 57 nsew signal output
rlabel metal2 s 6918 9840 6974 10000 6 N2BEGb[5]
port 58 nsew signal output
rlabel metal2 s 7286 9840 7342 10000 6 N2BEGb[6]
port 59 nsew signal output
rlabel metal2 s 7654 9840 7710 10000 6 N2BEGb[7]
port 60 nsew signal output
rlabel metal2 s 8022 9840 8078 10000 6 N4BEG[0]
port 61 nsew signal output
rlabel metal2 s 11702 9840 11758 10000 6 N4BEG[10]
port 62 nsew signal output
rlabel metal2 s 12070 9840 12126 10000 6 N4BEG[11]
port 63 nsew signal output
rlabel metal2 s 12438 9840 12494 10000 6 N4BEG[12]
port 64 nsew signal output
rlabel metal2 s 12806 9840 12862 10000 6 N4BEG[13]
port 65 nsew signal output
rlabel metal2 s 13174 9840 13230 10000 6 N4BEG[14]
port 66 nsew signal output
rlabel metal2 s 13542 9840 13598 10000 6 N4BEG[15]
port 67 nsew signal output
rlabel metal2 s 8390 9840 8446 10000 6 N4BEG[1]
port 68 nsew signal output
rlabel metal2 s 8758 9840 8814 10000 6 N4BEG[2]
port 69 nsew signal output
rlabel metal2 s 9126 9840 9182 10000 6 N4BEG[3]
port 70 nsew signal output
rlabel metal2 s 9494 9840 9550 10000 6 N4BEG[4]
port 71 nsew signal output
rlabel metal2 s 9862 9840 9918 10000 6 N4BEG[5]
port 72 nsew signal output
rlabel metal2 s 10230 9840 10286 10000 6 N4BEG[6]
port 73 nsew signal output
rlabel metal2 s 10598 9840 10654 10000 6 N4BEG[7]
port 74 nsew signal output
rlabel metal2 s 10966 9840 11022 10000 6 N4BEG[8]
port 75 nsew signal output
rlabel metal2 s 11334 9840 11390 10000 6 N4BEG[9]
port 76 nsew signal output
rlabel metal2 s 13910 9840 13966 10000 6 NN4BEG[0]
port 77 nsew signal output
rlabel metal2 s 17590 9840 17646 10000 6 NN4BEG[10]
port 78 nsew signal output
rlabel metal2 s 17958 9840 18014 10000 6 NN4BEG[11]
port 79 nsew signal output
rlabel metal2 s 18326 9840 18382 10000 6 NN4BEG[12]
port 80 nsew signal output
rlabel metal2 s 18694 9840 18750 10000 6 NN4BEG[13]
port 81 nsew signal output
rlabel metal2 s 19062 9840 19118 10000 6 NN4BEG[14]
port 82 nsew signal output
rlabel metal2 s 19430 9840 19486 10000 6 NN4BEG[15]
port 83 nsew signal output
rlabel metal2 s 14278 9840 14334 10000 6 NN4BEG[1]
port 84 nsew signal output
rlabel metal2 s 14646 9840 14702 10000 6 NN4BEG[2]
port 85 nsew signal output
rlabel metal2 s 15014 9840 15070 10000 6 NN4BEG[3]
port 86 nsew signal output
rlabel metal2 s 15382 9840 15438 10000 6 NN4BEG[4]
port 87 nsew signal output
rlabel metal2 s 15750 9840 15806 10000 6 NN4BEG[5]
port 88 nsew signal output
rlabel metal2 s 16118 9840 16174 10000 6 NN4BEG[6]
port 89 nsew signal output
rlabel metal2 s 16486 9840 16542 10000 6 NN4BEG[7]
port 90 nsew signal output
rlabel metal2 s 16854 9840 16910 10000 6 NN4BEG[8]
port 91 nsew signal output
rlabel metal2 s 17222 9840 17278 10000 6 NN4BEG[9]
port 92 nsew signal output
rlabel metal2 s 19798 9840 19854 10000 6 S1END[0]
port 93 nsew signal input
rlabel metal2 s 20166 9840 20222 10000 6 S1END[1]
port 94 nsew signal input
rlabel metal2 s 20534 9840 20590 10000 6 S1END[2]
port 95 nsew signal input
rlabel metal2 s 20902 9840 20958 10000 6 S1END[3]
port 96 nsew signal input
rlabel metal2 s 21270 9840 21326 10000 6 S2END[0]
port 97 nsew signal input
rlabel metal2 s 21638 9840 21694 10000 6 S2END[1]
port 98 nsew signal input
rlabel metal2 s 22006 9840 22062 10000 6 S2END[2]
port 99 nsew signal input
rlabel metal2 s 22374 9840 22430 10000 6 S2END[3]
port 100 nsew signal input
rlabel metal2 s 22742 9840 22798 10000 6 S2END[4]
port 101 nsew signal input
rlabel metal2 s 23110 9840 23166 10000 6 S2END[5]
port 102 nsew signal input
rlabel metal2 s 23478 9840 23534 10000 6 S2END[6]
port 103 nsew signal input
rlabel metal2 s 23846 9840 23902 10000 6 S2END[7]
port 104 nsew signal input
rlabel metal2 s 24214 9840 24270 10000 6 S2MID[0]
port 105 nsew signal input
rlabel metal2 s 24582 9840 24638 10000 6 S2MID[1]
port 106 nsew signal input
rlabel metal2 s 24950 9840 25006 10000 6 S2MID[2]
port 107 nsew signal input
rlabel metal2 s 25318 9840 25374 10000 6 S2MID[3]
port 108 nsew signal input
rlabel metal2 s 25686 9840 25742 10000 6 S2MID[4]
port 109 nsew signal input
rlabel metal2 s 26054 9840 26110 10000 6 S2MID[5]
port 110 nsew signal input
rlabel metal2 s 26422 9840 26478 10000 6 S2MID[6]
port 111 nsew signal input
rlabel metal2 s 26790 9840 26846 10000 6 S2MID[7]
port 112 nsew signal input
rlabel metal2 s 27158 9840 27214 10000 6 S4END[0]
port 113 nsew signal input
rlabel metal2 s 30838 9840 30894 10000 6 S4END[10]
port 114 nsew signal input
rlabel metal2 s 31206 9840 31262 10000 6 S4END[11]
port 115 nsew signal input
rlabel metal2 s 31574 9840 31630 10000 6 S4END[12]
port 116 nsew signal input
rlabel metal2 s 31942 9840 31998 10000 6 S4END[13]
port 117 nsew signal input
rlabel metal2 s 32310 9840 32366 10000 6 S4END[14]
port 118 nsew signal input
rlabel metal2 s 32678 9840 32734 10000 6 S4END[15]
port 119 nsew signal input
rlabel metal2 s 27526 9840 27582 10000 6 S4END[1]
port 120 nsew signal input
rlabel metal2 s 27894 9840 27950 10000 6 S4END[2]
port 121 nsew signal input
rlabel metal2 s 28262 9840 28318 10000 6 S4END[3]
port 122 nsew signal input
rlabel metal2 s 28630 9840 28686 10000 6 S4END[4]
port 123 nsew signal input
rlabel metal2 s 28998 9840 29054 10000 6 S4END[5]
port 124 nsew signal input
rlabel metal2 s 29366 9840 29422 10000 6 S4END[6]
port 125 nsew signal input
rlabel metal2 s 29734 9840 29790 10000 6 S4END[7]
port 126 nsew signal input
rlabel metal2 s 30102 9840 30158 10000 6 S4END[8]
port 127 nsew signal input
rlabel metal2 s 30470 9840 30526 10000 6 S4END[9]
port 128 nsew signal input
rlabel metal2 s 33046 9840 33102 10000 6 SS4END[0]
port 129 nsew signal input
rlabel metal2 s 36726 9840 36782 10000 6 SS4END[10]
port 130 nsew signal input
rlabel metal2 s 37094 9840 37150 10000 6 SS4END[11]
port 131 nsew signal input
rlabel metal2 s 37462 9840 37518 10000 6 SS4END[12]
port 132 nsew signal input
rlabel metal2 s 37830 9840 37886 10000 6 SS4END[13]
port 133 nsew signal input
rlabel metal2 s 38198 9840 38254 10000 6 SS4END[14]
port 134 nsew signal input
rlabel metal2 s 38566 9840 38622 10000 6 SS4END[15]
port 135 nsew signal input
rlabel metal2 s 33414 9840 33470 10000 6 SS4END[1]
port 136 nsew signal input
rlabel metal2 s 33782 9840 33838 10000 6 SS4END[2]
port 137 nsew signal input
rlabel metal2 s 34150 9840 34206 10000 6 SS4END[3]
port 138 nsew signal input
rlabel metal2 s 34518 9840 34574 10000 6 SS4END[4]
port 139 nsew signal input
rlabel metal2 s 34886 9840 34942 10000 6 SS4END[5]
port 140 nsew signal input
rlabel metal2 s 35254 9840 35310 10000 6 SS4END[6]
port 141 nsew signal input
rlabel metal2 s 35622 9840 35678 10000 6 SS4END[7]
port 142 nsew signal input
rlabel metal2 s 35990 9840 36046 10000 6 SS4END[8]
port 143 nsew signal input
rlabel metal2 s 36358 9840 36414 10000 6 SS4END[9]
port 144 nsew signal input
rlabel metal2 s 1398 0 1454 160 6 UserCLK
port 145 nsew signal input
rlabel metal2 s 38934 9840 38990 10000 6 UserCLKo
port 146 nsew signal output
rlabel metal4 s 6533 1040 6853 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 17711 1040 18031 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 28889 1040 29209 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 40067 1040 40387 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 12122 1040 12442 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 23300 1040 23620 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 34478 1040 34798 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 45656 1040 45976 8752 6 vssd1
port 148 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 47000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 584030
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/S_term_single2/runs/24_12_05_10_25/results/signoff/S_term_single2.magic.gds
string GDS_START 45964
<< end >>

