magic
tech sky130A
magscale 1 2
timestamp 1733394512
<< obsli1 >>
rect 1104 1071 45816 43537
<< obsm1 >>
rect 14 280 46998 43648
<< metal2 >>
rect 662 44840 718 45000
rect 1030 44840 1086 45000
rect 1398 44840 1454 45000
rect 1766 44840 1822 45000
rect 2134 44840 2190 45000
rect 2502 44840 2558 45000
rect 2870 44840 2926 45000
rect 3238 44840 3294 45000
rect 3606 44840 3662 45000
rect 3974 44840 4030 45000
rect 4342 44840 4398 45000
rect 4710 44840 4766 45000
rect 5078 44840 5134 45000
rect 5446 44840 5502 45000
rect 5814 44840 5870 45000
rect 6182 44840 6238 45000
rect 6550 44840 6606 45000
rect 6918 44840 6974 45000
rect 7286 44840 7342 45000
rect 7654 44840 7710 45000
rect 8022 44840 8078 45000
rect 8390 44840 8446 45000
rect 8758 44840 8814 45000
rect 9126 44840 9182 45000
rect 9494 44840 9550 45000
rect 9862 44840 9918 45000
rect 10230 44840 10286 45000
rect 10598 44840 10654 45000
rect 10966 44840 11022 45000
rect 11334 44840 11390 45000
rect 11702 44840 11758 45000
rect 12070 44840 12126 45000
rect 12438 44840 12494 45000
rect 12806 44840 12862 45000
rect 13174 44840 13230 45000
rect 13542 44840 13598 45000
rect 13910 44840 13966 45000
rect 14278 44840 14334 45000
rect 14646 44840 14702 45000
rect 15014 44840 15070 45000
rect 15382 44840 15438 45000
rect 15750 44840 15806 45000
rect 16118 44840 16174 45000
rect 16486 44840 16542 45000
rect 16854 44840 16910 45000
rect 17222 44840 17278 45000
rect 17590 44840 17646 45000
rect 17958 44840 18014 45000
rect 18326 44840 18382 45000
rect 18694 44840 18750 45000
rect 19062 44840 19118 45000
rect 19430 44840 19486 45000
rect 19798 44840 19854 45000
rect 20166 44840 20222 45000
rect 20534 44840 20590 45000
rect 20902 44840 20958 45000
rect 21270 44840 21326 45000
rect 21638 44840 21694 45000
rect 22006 44840 22062 45000
rect 22374 44840 22430 45000
rect 22742 44840 22798 45000
rect 23110 44840 23166 45000
rect 23478 44840 23534 45000
rect 23846 44840 23902 45000
rect 24214 44840 24270 45000
rect 24582 44840 24638 45000
rect 24950 44840 25006 45000
rect 25318 44840 25374 45000
rect 25686 44840 25742 45000
rect 26054 44840 26110 45000
rect 26422 44840 26478 45000
rect 26790 44840 26846 45000
rect 27158 44840 27214 45000
rect 27526 44840 27582 45000
rect 27894 44840 27950 45000
rect 28262 44840 28318 45000
rect 28630 44840 28686 45000
rect 28998 44840 29054 45000
rect 29366 44840 29422 45000
rect 29734 44840 29790 45000
rect 30102 44840 30158 45000
rect 30470 44840 30526 45000
rect 30838 44840 30894 45000
rect 31206 44840 31262 45000
rect 31574 44840 31630 45000
rect 31942 44840 31998 45000
rect 32310 44840 32366 45000
rect 32678 44840 32734 45000
rect 33046 44840 33102 45000
rect 33414 44840 33470 45000
rect 33782 44840 33838 45000
rect 34150 44840 34206 45000
rect 34518 44840 34574 45000
rect 34886 44840 34942 45000
rect 35254 44840 35310 45000
rect 35622 44840 35678 45000
rect 35990 44840 36046 45000
rect 36358 44840 36414 45000
rect 36726 44840 36782 45000
rect 37094 44840 37150 45000
rect 37462 44840 37518 45000
rect 37830 44840 37886 45000
rect 38198 44840 38254 45000
rect 38566 44840 38622 45000
rect 38934 44840 38990 45000
rect 39302 44840 39358 45000
rect 39670 44840 39726 45000
rect 40038 44840 40094 45000
rect 40406 44840 40462 45000
rect 40774 44840 40830 45000
rect 41142 44840 41198 45000
rect 41510 44840 41566 45000
rect 41878 44840 41934 45000
rect 42246 44840 42302 45000
rect 42614 44840 42670 45000
rect 42982 44840 43038 45000
rect 43350 44840 43406 45000
rect 43718 44840 43774 45000
rect 44086 44840 44142 45000
rect 44454 44840 44510 45000
rect 44822 44840 44878 45000
rect 45190 44840 45246 45000
rect 45558 44840 45614 45000
rect 45926 44840 45982 45000
rect 46294 44840 46350 45000
rect 662 0 718 160
rect 1030 0 1086 160
rect 1398 0 1454 160
rect 1766 0 1822 160
rect 2134 0 2190 160
rect 2502 0 2558 160
rect 2870 0 2926 160
rect 3238 0 3294 160
rect 3606 0 3662 160
rect 3974 0 4030 160
rect 4342 0 4398 160
rect 4710 0 4766 160
rect 5078 0 5134 160
rect 5446 0 5502 160
rect 5814 0 5870 160
rect 6182 0 6238 160
rect 6550 0 6606 160
rect 6918 0 6974 160
rect 7286 0 7342 160
rect 7654 0 7710 160
rect 8022 0 8078 160
rect 8390 0 8446 160
rect 8758 0 8814 160
rect 9126 0 9182 160
rect 9494 0 9550 160
rect 9862 0 9918 160
rect 10230 0 10286 160
rect 10598 0 10654 160
rect 10966 0 11022 160
rect 11334 0 11390 160
rect 11702 0 11758 160
rect 12070 0 12126 160
rect 12438 0 12494 160
rect 12806 0 12862 160
rect 13174 0 13230 160
rect 13542 0 13598 160
rect 13910 0 13966 160
rect 14278 0 14334 160
rect 14646 0 14702 160
rect 15014 0 15070 160
rect 15382 0 15438 160
rect 15750 0 15806 160
rect 16118 0 16174 160
rect 16486 0 16542 160
rect 16854 0 16910 160
rect 17222 0 17278 160
rect 17590 0 17646 160
rect 17958 0 18014 160
rect 18326 0 18382 160
rect 18694 0 18750 160
rect 19062 0 19118 160
rect 19430 0 19486 160
rect 19798 0 19854 160
rect 20166 0 20222 160
rect 20534 0 20590 160
rect 20902 0 20958 160
rect 21270 0 21326 160
rect 21638 0 21694 160
rect 22006 0 22062 160
rect 22374 0 22430 160
rect 22742 0 22798 160
rect 23110 0 23166 160
rect 23478 0 23534 160
rect 23846 0 23902 160
rect 24214 0 24270 160
rect 24582 0 24638 160
rect 24950 0 25006 160
rect 25318 0 25374 160
rect 25686 0 25742 160
rect 26054 0 26110 160
rect 26422 0 26478 160
rect 26790 0 26846 160
rect 27158 0 27214 160
rect 27526 0 27582 160
rect 27894 0 27950 160
rect 28262 0 28318 160
rect 28630 0 28686 160
rect 28998 0 29054 160
rect 29366 0 29422 160
rect 29734 0 29790 160
rect 30102 0 30158 160
rect 30470 0 30526 160
rect 30838 0 30894 160
rect 31206 0 31262 160
rect 31574 0 31630 160
rect 31942 0 31998 160
rect 32310 0 32366 160
rect 32678 0 32734 160
rect 33046 0 33102 160
rect 33414 0 33470 160
rect 33782 0 33838 160
rect 34150 0 34206 160
rect 34518 0 34574 160
rect 34886 0 34942 160
rect 35254 0 35310 160
rect 35622 0 35678 160
rect 35990 0 36046 160
rect 36358 0 36414 160
rect 36726 0 36782 160
rect 37094 0 37150 160
rect 37462 0 37518 160
rect 37830 0 37886 160
rect 38198 0 38254 160
rect 38566 0 38622 160
rect 38934 0 38990 160
rect 39302 0 39358 160
rect 39670 0 39726 160
rect 40038 0 40094 160
rect 40406 0 40462 160
rect 40774 0 40830 160
rect 41142 0 41198 160
rect 41510 0 41566 160
rect 41878 0 41934 160
rect 42246 0 42302 160
rect 42614 0 42670 160
rect 42982 0 43038 160
rect 43350 0 43406 160
rect 43718 0 43774 160
rect 44086 0 44142 160
rect 44454 0 44510 160
rect 44822 0 44878 160
rect 45190 0 45246 160
rect 45558 0 45614 160
rect 45926 0 45982 160
rect 46294 0 46350 160
<< obsm2 >>
rect 20 44784 606 44962
rect 774 44784 974 44962
rect 1142 44784 1342 44962
rect 1510 44784 1710 44962
rect 1878 44784 2078 44962
rect 2246 44784 2446 44962
rect 2614 44784 2814 44962
rect 2982 44784 3182 44962
rect 3350 44784 3550 44962
rect 3718 44784 3918 44962
rect 4086 44784 4286 44962
rect 4454 44784 4654 44962
rect 4822 44784 5022 44962
rect 5190 44784 5390 44962
rect 5558 44784 5758 44962
rect 5926 44784 6126 44962
rect 6294 44784 6494 44962
rect 6662 44784 6862 44962
rect 7030 44784 7230 44962
rect 7398 44784 7598 44962
rect 7766 44784 7966 44962
rect 8134 44784 8334 44962
rect 8502 44784 8702 44962
rect 8870 44784 9070 44962
rect 9238 44784 9438 44962
rect 9606 44784 9806 44962
rect 9974 44784 10174 44962
rect 10342 44784 10542 44962
rect 10710 44784 10910 44962
rect 11078 44784 11278 44962
rect 11446 44784 11646 44962
rect 11814 44784 12014 44962
rect 12182 44784 12382 44962
rect 12550 44784 12750 44962
rect 12918 44784 13118 44962
rect 13286 44784 13486 44962
rect 13654 44784 13854 44962
rect 14022 44784 14222 44962
rect 14390 44784 14590 44962
rect 14758 44784 14958 44962
rect 15126 44784 15326 44962
rect 15494 44784 15694 44962
rect 15862 44784 16062 44962
rect 16230 44784 16430 44962
rect 16598 44784 16798 44962
rect 16966 44784 17166 44962
rect 17334 44784 17534 44962
rect 17702 44784 17902 44962
rect 18070 44784 18270 44962
rect 18438 44784 18638 44962
rect 18806 44784 19006 44962
rect 19174 44784 19374 44962
rect 19542 44784 19742 44962
rect 19910 44784 20110 44962
rect 20278 44784 20478 44962
rect 20646 44784 20846 44962
rect 21014 44784 21214 44962
rect 21382 44784 21582 44962
rect 21750 44784 21950 44962
rect 22118 44784 22318 44962
rect 22486 44784 22686 44962
rect 22854 44784 23054 44962
rect 23222 44784 23422 44962
rect 23590 44784 23790 44962
rect 23958 44784 24158 44962
rect 24326 44784 24526 44962
rect 24694 44784 24894 44962
rect 25062 44784 25262 44962
rect 25430 44784 25630 44962
rect 25798 44784 25998 44962
rect 26166 44784 26366 44962
rect 26534 44784 26734 44962
rect 26902 44784 27102 44962
rect 27270 44784 27470 44962
rect 27638 44784 27838 44962
rect 28006 44784 28206 44962
rect 28374 44784 28574 44962
rect 28742 44784 28942 44962
rect 29110 44784 29310 44962
rect 29478 44784 29678 44962
rect 29846 44784 30046 44962
rect 30214 44784 30414 44962
rect 30582 44784 30782 44962
rect 30950 44784 31150 44962
rect 31318 44784 31518 44962
rect 31686 44784 31886 44962
rect 32054 44784 32254 44962
rect 32422 44784 32622 44962
rect 32790 44784 32990 44962
rect 33158 44784 33358 44962
rect 33526 44784 33726 44962
rect 33894 44784 34094 44962
rect 34262 44784 34462 44962
rect 34630 44784 34830 44962
rect 34998 44784 35198 44962
rect 35366 44784 35566 44962
rect 35734 44784 35934 44962
rect 36102 44784 36302 44962
rect 36470 44784 36670 44962
rect 36838 44784 37038 44962
rect 37206 44784 37406 44962
rect 37574 44784 37774 44962
rect 37942 44784 38142 44962
rect 38310 44784 38510 44962
rect 38678 44784 38878 44962
rect 39046 44784 39246 44962
rect 39414 44784 39614 44962
rect 39782 44784 39982 44962
rect 40150 44784 40350 44962
rect 40518 44784 40718 44962
rect 40886 44784 41086 44962
rect 41254 44784 41454 44962
rect 41622 44784 41822 44962
rect 41990 44784 42190 44962
rect 42358 44784 42558 44962
rect 42726 44784 42926 44962
rect 43094 44784 43294 44962
rect 43462 44784 43662 44962
rect 43830 44784 44030 44962
rect 44198 44784 44398 44962
rect 44566 44784 44766 44962
rect 44934 44784 45134 44962
rect 45302 44784 45502 44962
rect 45670 44784 45870 44962
rect 46038 44784 46238 44962
rect 46406 44784 46992 44962
rect 20 216 46992 44784
rect 20 54 606 216
rect 774 54 974 216
rect 1142 54 1342 216
rect 1510 54 1710 216
rect 1878 54 2078 216
rect 2246 54 2446 216
rect 2614 54 2814 216
rect 2982 54 3182 216
rect 3350 54 3550 216
rect 3718 54 3918 216
rect 4086 54 4286 216
rect 4454 54 4654 216
rect 4822 54 5022 216
rect 5190 54 5390 216
rect 5558 54 5758 216
rect 5926 54 6126 216
rect 6294 54 6494 216
rect 6662 54 6862 216
rect 7030 54 7230 216
rect 7398 54 7598 216
rect 7766 54 7966 216
rect 8134 54 8334 216
rect 8502 54 8702 216
rect 8870 54 9070 216
rect 9238 54 9438 216
rect 9606 54 9806 216
rect 9974 54 10174 216
rect 10342 54 10542 216
rect 10710 54 10910 216
rect 11078 54 11278 216
rect 11446 54 11646 216
rect 11814 54 12014 216
rect 12182 54 12382 216
rect 12550 54 12750 216
rect 12918 54 13118 216
rect 13286 54 13486 216
rect 13654 54 13854 216
rect 14022 54 14222 216
rect 14390 54 14590 216
rect 14758 54 14958 216
rect 15126 54 15326 216
rect 15494 54 15694 216
rect 15862 54 16062 216
rect 16230 54 16430 216
rect 16598 54 16798 216
rect 16966 54 17166 216
rect 17334 54 17534 216
rect 17702 54 17902 216
rect 18070 54 18270 216
rect 18438 54 18638 216
rect 18806 54 19006 216
rect 19174 54 19374 216
rect 19542 54 19742 216
rect 19910 54 20110 216
rect 20278 54 20478 216
rect 20646 54 20846 216
rect 21014 54 21214 216
rect 21382 54 21582 216
rect 21750 54 21950 216
rect 22118 54 22318 216
rect 22486 54 22686 216
rect 22854 54 23054 216
rect 23222 54 23422 216
rect 23590 54 23790 216
rect 23958 54 24158 216
rect 24326 54 24526 216
rect 24694 54 24894 216
rect 25062 54 25262 216
rect 25430 54 25630 216
rect 25798 54 25998 216
rect 26166 54 26366 216
rect 26534 54 26734 216
rect 26902 54 27102 216
rect 27270 54 27470 216
rect 27638 54 27838 216
rect 28006 54 28206 216
rect 28374 54 28574 216
rect 28742 54 28942 216
rect 29110 54 29310 216
rect 29478 54 29678 216
rect 29846 54 30046 216
rect 30214 54 30414 216
rect 30582 54 30782 216
rect 30950 54 31150 216
rect 31318 54 31518 216
rect 31686 54 31886 216
rect 32054 54 32254 216
rect 32422 54 32622 216
rect 32790 54 32990 216
rect 33158 54 33358 216
rect 33526 54 33726 216
rect 33894 54 34094 216
rect 34262 54 34462 216
rect 34630 54 34830 216
rect 34998 54 35198 216
rect 35366 54 35566 216
rect 35734 54 35934 216
rect 36102 54 36302 216
rect 36470 54 36670 216
rect 36838 54 37038 216
rect 37206 54 37406 216
rect 37574 54 37774 216
rect 37942 54 38142 216
rect 38310 54 38510 216
rect 38678 54 38878 216
rect 39046 54 39246 216
rect 39414 54 39614 216
rect 39782 54 39982 216
rect 40150 54 40350 216
rect 40518 54 40718 216
rect 40886 54 41086 216
rect 41254 54 41454 216
rect 41622 54 41822 216
rect 41990 54 42190 216
rect 42358 54 42558 216
rect 42726 54 42926 216
rect 43094 54 43294 216
rect 43462 54 43662 216
rect 43830 54 44030 216
rect 44198 54 44398 216
rect 44566 54 44766 216
rect 44934 54 45134 216
rect 45302 54 45502 216
rect 45670 54 45870 216
rect 46038 54 46238 216
rect 46406 54 46992 216
<< metal3 >>
rect 0 39720 160 39840
rect 0 39448 160 39568
rect 0 39176 160 39296
rect 0 38904 160 39024
rect 0 38632 160 38752
rect 0 38360 160 38480
rect 0 38088 160 38208
rect 0 37816 160 37936
rect 0 37544 160 37664
rect 0 37272 160 37392
rect 0 37000 160 37120
rect 0 36728 160 36848
rect 0 36456 160 36576
rect 0 36184 160 36304
rect 0 35912 160 36032
rect 0 35640 160 35760
rect 0 35368 160 35488
rect 0 35096 160 35216
rect 0 34824 160 34944
rect 0 34552 160 34672
rect 0 34280 160 34400
rect 0 34008 160 34128
rect 0 33736 160 33856
rect 0 33464 160 33584
rect 0 33192 160 33312
rect 0 32920 160 33040
rect 0 32648 160 32768
rect 0 32376 160 32496
rect 0 32104 160 32224
rect 0 31832 160 31952
rect 0 31560 160 31680
rect 0 31288 160 31408
rect 0 31016 160 31136
rect 0 30744 160 30864
rect 0 30472 160 30592
rect 0 30200 160 30320
rect 0 29928 160 30048
rect 0 29656 160 29776
rect 0 29384 160 29504
rect 0 29112 160 29232
rect 0 28840 160 28960
rect 0 28568 160 28688
rect 0 28296 160 28416
rect 0 28024 160 28144
rect 0 27752 160 27872
rect 0 27480 160 27600
rect 0 27208 160 27328
rect 0 26936 160 27056
rect 0 26664 160 26784
rect 0 26392 160 26512
rect 0 26120 160 26240
rect 0 25848 160 25968
rect 0 25576 160 25696
rect 0 25304 160 25424
rect 0 25032 160 25152
rect 0 24760 160 24880
rect 0 24488 160 24608
rect 0 24216 160 24336
rect 0 23944 160 24064
rect 0 23672 160 23792
rect 0 23400 160 23520
rect 0 23128 160 23248
rect 0 22856 160 22976
rect 0 22584 160 22704
rect 0 22312 160 22432
rect 0 22040 160 22160
rect 0 21768 160 21888
rect 0 21496 160 21616
rect 0 21224 160 21344
rect 0 20952 160 21072
rect 0 20680 160 20800
rect 0 20408 160 20528
rect 0 20136 160 20256
rect 0 19864 160 19984
rect 0 19592 160 19712
rect 0 19320 160 19440
rect 0 19048 160 19168
rect 0 18776 160 18896
rect 0 18504 160 18624
rect 0 18232 160 18352
rect 0 17960 160 18080
rect 0 17688 160 17808
rect 0 17416 160 17536
rect 0 17144 160 17264
rect 0 16872 160 16992
rect 0 16600 160 16720
rect 0 16328 160 16448
rect 0 16056 160 16176
rect 0 15784 160 15904
rect 0 15512 160 15632
rect 0 15240 160 15360
rect 0 14968 160 15088
rect 0 14696 160 14816
rect 0 14424 160 14544
rect 0 14152 160 14272
rect 0 13880 160 14000
rect 0 13608 160 13728
rect 0 13336 160 13456
rect 0 13064 160 13184
rect 0 12792 160 12912
rect 0 12520 160 12640
rect 0 12248 160 12368
rect 0 11976 160 12096
rect 0 11704 160 11824
rect 0 11432 160 11552
rect 0 11160 160 11280
rect 0 10888 160 11008
rect 0 10616 160 10736
rect 0 10344 160 10464
rect 0 10072 160 10192
rect 0 9800 160 9920
rect 0 9528 160 9648
rect 0 9256 160 9376
rect 0 8984 160 9104
rect 0 8712 160 8832
rect 0 8440 160 8560
rect 0 8168 160 8288
rect 0 7896 160 8016
rect 0 7624 160 7744
rect 0 7352 160 7472
rect 0 7080 160 7200
rect 0 6808 160 6928
rect 0 6536 160 6656
rect 0 6264 160 6384
rect 0 5992 160 6112
rect 0 5720 160 5840
rect 0 5448 160 5568
rect 0 5176 160 5296
rect 46840 39720 47000 39840
rect 46840 39448 47000 39568
rect 46840 39176 47000 39296
rect 46840 38904 47000 39024
rect 46840 38632 47000 38752
rect 46840 38360 47000 38480
rect 46840 38088 47000 38208
rect 46840 37816 47000 37936
rect 46840 37544 47000 37664
rect 46840 37272 47000 37392
rect 46840 37000 47000 37120
rect 46840 36728 47000 36848
rect 46840 36456 47000 36576
rect 46840 36184 47000 36304
rect 46840 35912 47000 36032
rect 46840 35640 47000 35760
rect 46840 35368 47000 35488
rect 46840 35096 47000 35216
rect 46840 34824 47000 34944
rect 46840 34552 47000 34672
rect 46840 34280 47000 34400
rect 46840 34008 47000 34128
rect 46840 33736 47000 33856
rect 46840 33464 47000 33584
rect 46840 33192 47000 33312
rect 46840 32920 47000 33040
rect 46840 32648 47000 32768
rect 46840 32376 47000 32496
rect 46840 32104 47000 32224
rect 46840 31832 47000 31952
rect 46840 31560 47000 31680
rect 46840 31288 47000 31408
rect 46840 31016 47000 31136
rect 46840 30744 47000 30864
rect 46840 30472 47000 30592
rect 46840 30200 47000 30320
rect 46840 29928 47000 30048
rect 46840 29656 47000 29776
rect 46840 29384 47000 29504
rect 46840 29112 47000 29232
rect 46840 28840 47000 28960
rect 46840 28568 47000 28688
rect 46840 28296 47000 28416
rect 46840 28024 47000 28144
rect 46840 27752 47000 27872
rect 46840 27480 47000 27600
rect 46840 27208 47000 27328
rect 46840 26936 47000 27056
rect 46840 26664 47000 26784
rect 46840 26392 47000 26512
rect 46840 26120 47000 26240
rect 46840 25848 47000 25968
rect 46840 25576 47000 25696
rect 46840 25304 47000 25424
rect 46840 25032 47000 25152
rect 46840 24760 47000 24880
rect 46840 24488 47000 24608
rect 46840 24216 47000 24336
rect 46840 23944 47000 24064
rect 46840 23672 47000 23792
rect 46840 23400 47000 23520
rect 46840 23128 47000 23248
rect 46840 22856 47000 22976
rect 46840 22584 47000 22704
rect 46840 22312 47000 22432
rect 46840 22040 47000 22160
rect 46840 21768 47000 21888
rect 46840 21496 47000 21616
rect 46840 21224 47000 21344
rect 46840 20952 47000 21072
rect 46840 20680 47000 20800
rect 46840 20408 47000 20528
rect 46840 20136 47000 20256
rect 46840 19864 47000 19984
rect 46840 19592 47000 19712
rect 46840 19320 47000 19440
rect 46840 19048 47000 19168
rect 46840 18776 47000 18896
rect 46840 18504 47000 18624
rect 46840 18232 47000 18352
rect 46840 17960 47000 18080
rect 46840 17688 47000 17808
rect 46840 17416 47000 17536
rect 46840 17144 47000 17264
rect 46840 16872 47000 16992
rect 46840 16600 47000 16720
rect 46840 16328 47000 16448
rect 46840 16056 47000 16176
rect 46840 15784 47000 15904
rect 46840 15512 47000 15632
rect 46840 15240 47000 15360
rect 46840 14968 47000 15088
rect 46840 14696 47000 14816
rect 46840 14424 47000 14544
rect 46840 14152 47000 14272
rect 46840 13880 47000 14000
rect 46840 13608 47000 13728
rect 46840 13336 47000 13456
rect 46840 13064 47000 13184
rect 46840 12792 47000 12912
rect 46840 12520 47000 12640
rect 46840 12248 47000 12368
rect 46840 11976 47000 12096
rect 46840 11704 47000 11824
rect 46840 11432 47000 11552
rect 46840 11160 47000 11280
rect 46840 10888 47000 11008
rect 46840 10616 47000 10736
rect 46840 10344 47000 10464
rect 46840 10072 47000 10192
rect 46840 9800 47000 9920
rect 46840 9528 47000 9648
rect 46840 9256 47000 9376
rect 46840 8984 47000 9104
rect 46840 8712 47000 8832
rect 46840 8440 47000 8560
rect 46840 8168 47000 8288
rect 46840 7896 47000 8016
rect 46840 7624 47000 7744
rect 46840 7352 47000 7472
rect 46840 7080 47000 7200
rect 46840 6808 47000 6928
rect 46840 6536 47000 6656
rect 46840 6264 47000 6384
rect 46840 5992 47000 6112
rect 46840 5720 47000 5840
rect 46840 5448 47000 5568
rect 46840 5176 47000 5296
<< obsm3 >>
rect 160 39920 46907 43553
rect 240 5096 46760 39920
rect 160 1055 46907 5096
<< metal4 >>
rect 4208 1040 4528 43568
rect 19568 1040 19888 43568
rect 34928 1040 35248 43568
<< obsm4 >>
rect 427 1123 4128 43213
rect 4608 1123 19488 43213
rect 19968 1123 34848 43213
rect 35328 1123 46309 43213
<< labels >>
rlabel metal3 s 46840 18232 47000 18352 6 E1BEG[0]
port 1 nsew signal output
rlabel metal3 s 46840 18504 47000 18624 6 E1BEG[1]
port 2 nsew signal output
rlabel metal3 s 46840 18776 47000 18896 6 E1BEG[2]
port 3 nsew signal output
rlabel metal3 s 46840 19048 47000 19168 6 E1BEG[3]
port 4 nsew signal output
rlabel metal3 s 0 18232 160 18352 6 E1END[0]
port 5 nsew signal input
rlabel metal3 s 0 18504 160 18624 6 E1END[1]
port 6 nsew signal input
rlabel metal3 s 0 18776 160 18896 6 E1END[2]
port 7 nsew signal input
rlabel metal3 s 0 19048 160 19168 6 E1END[3]
port 8 nsew signal input
rlabel metal3 s 46840 19320 47000 19440 6 E2BEG[0]
port 9 nsew signal output
rlabel metal3 s 46840 19592 47000 19712 6 E2BEG[1]
port 10 nsew signal output
rlabel metal3 s 46840 19864 47000 19984 6 E2BEG[2]
port 11 nsew signal output
rlabel metal3 s 46840 20136 47000 20256 6 E2BEG[3]
port 12 nsew signal output
rlabel metal3 s 46840 20408 47000 20528 6 E2BEG[4]
port 13 nsew signal output
rlabel metal3 s 46840 20680 47000 20800 6 E2BEG[5]
port 14 nsew signal output
rlabel metal3 s 46840 20952 47000 21072 6 E2BEG[6]
port 15 nsew signal output
rlabel metal3 s 46840 21224 47000 21344 6 E2BEG[7]
port 16 nsew signal output
rlabel metal3 s 46840 21496 47000 21616 6 E2BEGb[0]
port 17 nsew signal output
rlabel metal3 s 46840 21768 47000 21888 6 E2BEGb[1]
port 18 nsew signal output
rlabel metal3 s 46840 22040 47000 22160 6 E2BEGb[2]
port 19 nsew signal output
rlabel metal3 s 46840 22312 47000 22432 6 E2BEGb[3]
port 20 nsew signal output
rlabel metal3 s 46840 22584 47000 22704 6 E2BEGb[4]
port 21 nsew signal output
rlabel metal3 s 46840 22856 47000 22976 6 E2BEGb[5]
port 22 nsew signal output
rlabel metal3 s 46840 23128 47000 23248 6 E2BEGb[6]
port 23 nsew signal output
rlabel metal3 s 46840 23400 47000 23520 6 E2BEGb[7]
port 24 nsew signal output
rlabel metal3 s 0 21496 160 21616 6 E2END[0]
port 25 nsew signal input
rlabel metal3 s 0 21768 160 21888 6 E2END[1]
port 26 nsew signal input
rlabel metal3 s 0 22040 160 22160 6 E2END[2]
port 27 nsew signal input
rlabel metal3 s 0 22312 160 22432 6 E2END[3]
port 28 nsew signal input
rlabel metal3 s 0 22584 160 22704 6 E2END[4]
port 29 nsew signal input
rlabel metal3 s 0 22856 160 22976 6 E2END[5]
port 30 nsew signal input
rlabel metal3 s 0 23128 160 23248 6 E2END[6]
port 31 nsew signal input
rlabel metal3 s 0 23400 160 23520 6 E2END[7]
port 32 nsew signal input
rlabel metal3 s 0 19320 160 19440 6 E2MID[0]
port 33 nsew signal input
rlabel metal3 s 0 19592 160 19712 6 E2MID[1]
port 34 nsew signal input
rlabel metal3 s 0 19864 160 19984 6 E2MID[2]
port 35 nsew signal input
rlabel metal3 s 0 20136 160 20256 6 E2MID[3]
port 36 nsew signal input
rlabel metal3 s 0 20408 160 20528 6 E2MID[4]
port 37 nsew signal input
rlabel metal3 s 0 20680 160 20800 6 E2MID[5]
port 38 nsew signal input
rlabel metal3 s 0 20952 160 21072 6 E2MID[6]
port 39 nsew signal input
rlabel metal3 s 0 21224 160 21344 6 E2MID[7]
port 40 nsew signal input
rlabel metal3 s 46840 28024 47000 28144 6 E6BEG[0]
port 41 nsew signal output
rlabel metal3 s 46840 30744 47000 30864 6 E6BEG[10]
port 42 nsew signal output
rlabel metal3 s 46840 31016 47000 31136 6 E6BEG[11]
port 43 nsew signal output
rlabel metal3 s 46840 28296 47000 28416 6 E6BEG[1]
port 44 nsew signal output
rlabel metal3 s 46840 28568 47000 28688 6 E6BEG[2]
port 45 nsew signal output
rlabel metal3 s 46840 28840 47000 28960 6 E6BEG[3]
port 46 nsew signal output
rlabel metal3 s 46840 29112 47000 29232 6 E6BEG[4]
port 47 nsew signal output
rlabel metal3 s 46840 29384 47000 29504 6 E6BEG[5]
port 48 nsew signal output
rlabel metal3 s 46840 29656 47000 29776 6 E6BEG[6]
port 49 nsew signal output
rlabel metal3 s 46840 29928 47000 30048 6 E6BEG[7]
port 50 nsew signal output
rlabel metal3 s 46840 30200 47000 30320 6 E6BEG[8]
port 51 nsew signal output
rlabel metal3 s 46840 30472 47000 30592 6 E6BEG[9]
port 52 nsew signal output
rlabel metal3 s 0 28024 160 28144 6 E6END[0]
port 53 nsew signal input
rlabel metal3 s 0 30744 160 30864 6 E6END[10]
port 54 nsew signal input
rlabel metal3 s 0 31016 160 31136 6 E6END[11]
port 55 nsew signal input
rlabel metal3 s 0 28296 160 28416 6 E6END[1]
port 56 nsew signal input
rlabel metal3 s 0 28568 160 28688 6 E6END[2]
port 57 nsew signal input
rlabel metal3 s 0 28840 160 28960 6 E6END[3]
port 58 nsew signal input
rlabel metal3 s 0 29112 160 29232 6 E6END[4]
port 59 nsew signal input
rlabel metal3 s 0 29384 160 29504 6 E6END[5]
port 60 nsew signal input
rlabel metal3 s 0 29656 160 29776 6 E6END[6]
port 61 nsew signal input
rlabel metal3 s 0 29928 160 30048 6 E6END[7]
port 62 nsew signal input
rlabel metal3 s 0 30200 160 30320 6 E6END[8]
port 63 nsew signal input
rlabel metal3 s 0 30472 160 30592 6 E6END[9]
port 64 nsew signal input
rlabel metal3 s 46840 23672 47000 23792 6 EE4BEG[0]
port 65 nsew signal output
rlabel metal3 s 46840 26392 47000 26512 6 EE4BEG[10]
port 66 nsew signal output
rlabel metal3 s 46840 26664 47000 26784 6 EE4BEG[11]
port 67 nsew signal output
rlabel metal3 s 46840 26936 47000 27056 6 EE4BEG[12]
port 68 nsew signal output
rlabel metal3 s 46840 27208 47000 27328 6 EE4BEG[13]
port 69 nsew signal output
rlabel metal3 s 46840 27480 47000 27600 6 EE4BEG[14]
port 70 nsew signal output
rlabel metal3 s 46840 27752 47000 27872 6 EE4BEG[15]
port 71 nsew signal output
rlabel metal3 s 46840 23944 47000 24064 6 EE4BEG[1]
port 72 nsew signal output
rlabel metal3 s 46840 24216 47000 24336 6 EE4BEG[2]
port 73 nsew signal output
rlabel metal3 s 46840 24488 47000 24608 6 EE4BEG[3]
port 74 nsew signal output
rlabel metal3 s 46840 24760 47000 24880 6 EE4BEG[4]
port 75 nsew signal output
rlabel metal3 s 46840 25032 47000 25152 6 EE4BEG[5]
port 76 nsew signal output
rlabel metal3 s 46840 25304 47000 25424 6 EE4BEG[6]
port 77 nsew signal output
rlabel metal3 s 46840 25576 47000 25696 6 EE4BEG[7]
port 78 nsew signal output
rlabel metal3 s 46840 25848 47000 25968 6 EE4BEG[8]
port 79 nsew signal output
rlabel metal3 s 46840 26120 47000 26240 6 EE4BEG[9]
port 80 nsew signal output
rlabel metal3 s 0 23672 160 23792 6 EE4END[0]
port 81 nsew signal input
rlabel metal3 s 0 26392 160 26512 6 EE4END[10]
port 82 nsew signal input
rlabel metal3 s 0 26664 160 26784 6 EE4END[11]
port 83 nsew signal input
rlabel metal3 s 0 26936 160 27056 6 EE4END[12]
port 84 nsew signal input
rlabel metal3 s 0 27208 160 27328 6 EE4END[13]
port 85 nsew signal input
rlabel metal3 s 0 27480 160 27600 6 EE4END[14]
port 86 nsew signal input
rlabel metal3 s 0 27752 160 27872 6 EE4END[15]
port 87 nsew signal input
rlabel metal3 s 0 23944 160 24064 6 EE4END[1]
port 88 nsew signal input
rlabel metal3 s 0 24216 160 24336 6 EE4END[2]
port 89 nsew signal input
rlabel metal3 s 0 24488 160 24608 6 EE4END[3]
port 90 nsew signal input
rlabel metal3 s 0 24760 160 24880 6 EE4END[4]
port 91 nsew signal input
rlabel metal3 s 0 25032 160 25152 6 EE4END[5]
port 92 nsew signal input
rlabel metal3 s 0 25304 160 25424 6 EE4END[6]
port 93 nsew signal input
rlabel metal3 s 0 25576 160 25696 6 EE4END[7]
port 94 nsew signal input
rlabel metal3 s 0 25848 160 25968 6 EE4END[8]
port 95 nsew signal input
rlabel metal3 s 0 26120 160 26240 6 EE4END[9]
port 96 nsew signal input
rlabel metal3 s 0 31288 160 31408 6 FrameData[0]
port 97 nsew signal input
rlabel metal3 s 0 34008 160 34128 6 FrameData[10]
port 98 nsew signal input
rlabel metal3 s 0 34280 160 34400 6 FrameData[11]
port 99 nsew signal input
rlabel metal3 s 0 34552 160 34672 6 FrameData[12]
port 100 nsew signal input
rlabel metal3 s 0 34824 160 34944 6 FrameData[13]
port 101 nsew signal input
rlabel metal3 s 0 35096 160 35216 6 FrameData[14]
port 102 nsew signal input
rlabel metal3 s 0 35368 160 35488 6 FrameData[15]
port 103 nsew signal input
rlabel metal3 s 0 35640 160 35760 6 FrameData[16]
port 104 nsew signal input
rlabel metal3 s 0 35912 160 36032 6 FrameData[17]
port 105 nsew signal input
rlabel metal3 s 0 36184 160 36304 6 FrameData[18]
port 106 nsew signal input
rlabel metal3 s 0 36456 160 36576 6 FrameData[19]
port 107 nsew signal input
rlabel metal3 s 0 31560 160 31680 6 FrameData[1]
port 108 nsew signal input
rlabel metal3 s 0 36728 160 36848 6 FrameData[20]
port 109 nsew signal input
rlabel metal3 s 0 37000 160 37120 6 FrameData[21]
port 110 nsew signal input
rlabel metal3 s 0 37272 160 37392 6 FrameData[22]
port 111 nsew signal input
rlabel metal3 s 0 37544 160 37664 6 FrameData[23]
port 112 nsew signal input
rlabel metal3 s 0 37816 160 37936 6 FrameData[24]
port 113 nsew signal input
rlabel metal3 s 0 38088 160 38208 6 FrameData[25]
port 114 nsew signal input
rlabel metal3 s 0 38360 160 38480 6 FrameData[26]
port 115 nsew signal input
rlabel metal3 s 0 38632 160 38752 6 FrameData[27]
port 116 nsew signal input
rlabel metal3 s 0 38904 160 39024 6 FrameData[28]
port 117 nsew signal input
rlabel metal3 s 0 39176 160 39296 6 FrameData[29]
port 118 nsew signal input
rlabel metal3 s 0 31832 160 31952 6 FrameData[2]
port 119 nsew signal input
rlabel metal3 s 0 39448 160 39568 6 FrameData[30]
port 120 nsew signal input
rlabel metal3 s 0 39720 160 39840 6 FrameData[31]
port 121 nsew signal input
rlabel metal3 s 0 32104 160 32224 6 FrameData[3]
port 122 nsew signal input
rlabel metal3 s 0 32376 160 32496 6 FrameData[4]
port 123 nsew signal input
rlabel metal3 s 0 32648 160 32768 6 FrameData[5]
port 124 nsew signal input
rlabel metal3 s 0 32920 160 33040 6 FrameData[6]
port 125 nsew signal input
rlabel metal3 s 0 33192 160 33312 6 FrameData[7]
port 126 nsew signal input
rlabel metal3 s 0 33464 160 33584 6 FrameData[8]
port 127 nsew signal input
rlabel metal3 s 0 33736 160 33856 6 FrameData[9]
port 128 nsew signal input
rlabel metal3 s 46840 31288 47000 31408 6 FrameData_O[0]
port 129 nsew signal output
rlabel metal3 s 46840 34008 47000 34128 6 FrameData_O[10]
port 130 nsew signal output
rlabel metal3 s 46840 34280 47000 34400 6 FrameData_O[11]
port 131 nsew signal output
rlabel metal3 s 46840 34552 47000 34672 6 FrameData_O[12]
port 132 nsew signal output
rlabel metal3 s 46840 34824 47000 34944 6 FrameData_O[13]
port 133 nsew signal output
rlabel metal3 s 46840 35096 47000 35216 6 FrameData_O[14]
port 134 nsew signal output
rlabel metal3 s 46840 35368 47000 35488 6 FrameData_O[15]
port 135 nsew signal output
rlabel metal3 s 46840 35640 47000 35760 6 FrameData_O[16]
port 136 nsew signal output
rlabel metal3 s 46840 35912 47000 36032 6 FrameData_O[17]
port 137 nsew signal output
rlabel metal3 s 46840 36184 47000 36304 6 FrameData_O[18]
port 138 nsew signal output
rlabel metal3 s 46840 36456 47000 36576 6 FrameData_O[19]
port 139 nsew signal output
rlabel metal3 s 46840 31560 47000 31680 6 FrameData_O[1]
port 140 nsew signal output
rlabel metal3 s 46840 36728 47000 36848 6 FrameData_O[20]
port 141 nsew signal output
rlabel metal3 s 46840 37000 47000 37120 6 FrameData_O[21]
port 142 nsew signal output
rlabel metal3 s 46840 37272 47000 37392 6 FrameData_O[22]
port 143 nsew signal output
rlabel metal3 s 46840 37544 47000 37664 6 FrameData_O[23]
port 144 nsew signal output
rlabel metal3 s 46840 37816 47000 37936 6 FrameData_O[24]
port 145 nsew signal output
rlabel metal3 s 46840 38088 47000 38208 6 FrameData_O[25]
port 146 nsew signal output
rlabel metal3 s 46840 38360 47000 38480 6 FrameData_O[26]
port 147 nsew signal output
rlabel metal3 s 46840 38632 47000 38752 6 FrameData_O[27]
port 148 nsew signal output
rlabel metal3 s 46840 38904 47000 39024 6 FrameData_O[28]
port 149 nsew signal output
rlabel metal3 s 46840 39176 47000 39296 6 FrameData_O[29]
port 150 nsew signal output
rlabel metal3 s 46840 31832 47000 31952 6 FrameData_O[2]
port 151 nsew signal output
rlabel metal3 s 46840 39448 47000 39568 6 FrameData_O[30]
port 152 nsew signal output
rlabel metal3 s 46840 39720 47000 39840 6 FrameData_O[31]
port 153 nsew signal output
rlabel metal3 s 46840 32104 47000 32224 6 FrameData_O[3]
port 154 nsew signal output
rlabel metal3 s 46840 32376 47000 32496 6 FrameData_O[4]
port 155 nsew signal output
rlabel metal3 s 46840 32648 47000 32768 6 FrameData_O[5]
port 156 nsew signal output
rlabel metal3 s 46840 32920 47000 33040 6 FrameData_O[6]
port 157 nsew signal output
rlabel metal3 s 46840 33192 47000 33312 6 FrameData_O[7]
port 158 nsew signal output
rlabel metal3 s 46840 33464 47000 33584 6 FrameData_O[8]
port 159 nsew signal output
rlabel metal3 s 46840 33736 47000 33856 6 FrameData_O[9]
port 160 nsew signal output
rlabel metal2 s 39302 0 39358 160 6 FrameStrobe[0]
port 161 nsew signal input
rlabel metal2 s 42982 0 43038 160 6 FrameStrobe[10]
port 162 nsew signal input
rlabel metal2 s 43350 0 43406 160 6 FrameStrobe[11]
port 163 nsew signal input
rlabel metal2 s 43718 0 43774 160 6 FrameStrobe[12]
port 164 nsew signal input
rlabel metal2 s 44086 0 44142 160 6 FrameStrobe[13]
port 165 nsew signal input
rlabel metal2 s 44454 0 44510 160 6 FrameStrobe[14]
port 166 nsew signal input
rlabel metal2 s 44822 0 44878 160 6 FrameStrobe[15]
port 167 nsew signal input
rlabel metal2 s 45190 0 45246 160 6 FrameStrobe[16]
port 168 nsew signal input
rlabel metal2 s 45558 0 45614 160 6 FrameStrobe[17]
port 169 nsew signal input
rlabel metal2 s 45926 0 45982 160 6 FrameStrobe[18]
port 170 nsew signal input
rlabel metal2 s 46294 0 46350 160 6 FrameStrobe[19]
port 171 nsew signal input
rlabel metal2 s 39670 0 39726 160 6 FrameStrobe[1]
port 172 nsew signal input
rlabel metal2 s 40038 0 40094 160 6 FrameStrobe[2]
port 173 nsew signal input
rlabel metal2 s 40406 0 40462 160 6 FrameStrobe[3]
port 174 nsew signal input
rlabel metal2 s 40774 0 40830 160 6 FrameStrobe[4]
port 175 nsew signal input
rlabel metal2 s 41142 0 41198 160 6 FrameStrobe[5]
port 176 nsew signal input
rlabel metal2 s 41510 0 41566 160 6 FrameStrobe[6]
port 177 nsew signal input
rlabel metal2 s 41878 0 41934 160 6 FrameStrobe[7]
port 178 nsew signal input
rlabel metal2 s 42246 0 42302 160 6 FrameStrobe[8]
port 179 nsew signal input
rlabel metal2 s 42614 0 42670 160 6 FrameStrobe[9]
port 180 nsew signal input
rlabel metal2 s 39302 44840 39358 45000 6 FrameStrobe_O[0]
port 181 nsew signal output
rlabel metal2 s 42982 44840 43038 45000 6 FrameStrobe_O[10]
port 182 nsew signal output
rlabel metal2 s 43350 44840 43406 45000 6 FrameStrobe_O[11]
port 183 nsew signal output
rlabel metal2 s 43718 44840 43774 45000 6 FrameStrobe_O[12]
port 184 nsew signal output
rlabel metal2 s 44086 44840 44142 45000 6 FrameStrobe_O[13]
port 185 nsew signal output
rlabel metal2 s 44454 44840 44510 45000 6 FrameStrobe_O[14]
port 186 nsew signal output
rlabel metal2 s 44822 44840 44878 45000 6 FrameStrobe_O[15]
port 187 nsew signal output
rlabel metal2 s 45190 44840 45246 45000 6 FrameStrobe_O[16]
port 188 nsew signal output
rlabel metal2 s 45558 44840 45614 45000 6 FrameStrobe_O[17]
port 189 nsew signal output
rlabel metal2 s 45926 44840 45982 45000 6 FrameStrobe_O[18]
port 190 nsew signal output
rlabel metal2 s 46294 44840 46350 45000 6 FrameStrobe_O[19]
port 191 nsew signal output
rlabel metal2 s 39670 44840 39726 45000 6 FrameStrobe_O[1]
port 192 nsew signal output
rlabel metal2 s 40038 44840 40094 45000 6 FrameStrobe_O[2]
port 193 nsew signal output
rlabel metal2 s 40406 44840 40462 45000 6 FrameStrobe_O[3]
port 194 nsew signal output
rlabel metal2 s 40774 44840 40830 45000 6 FrameStrobe_O[4]
port 195 nsew signal output
rlabel metal2 s 41142 44840 41198 45000 6 FrameStrobe_O[5]
port 196 nsew signal output
rlabel metal2 s 41510 44840 41566 45000 6 FrameStrobe_O[6]
port 197 nsew signal output
rlabel metal2 s 41878 44840 41934 45000 6 FrameStrobe_O[7]
port 198 nsew signal output
rlabel metal2 s 42246 44840 42302 45000 6 FrameStrobe_O[8]
port 199 nsew signal output
rlabel metal2 s 42614 44840 42670 45000 6 FrameStrobe_O[9]
port 200 nsew signal output
rlabel metal2 s 662 44840 718 45000 6 N1BEG[0]
port 201 nsew signal output
rlabel metal2 s 1030 44840 1086 45000 6 N1BEG[1]
port 202 nsew signal output
rlabel metal2 s 1398 44840 1454 45000 6 N1BEG[2]
port 203 nsew signal output
rlabel metal2 s 1766 44840 1822 45000 6 N1BEG[3]
port 204 nsew signal output
rlabel metal2 s 662 0 718 160 6 N1END[0]
port 205 nsew signal input
rlabel metal2 s 1030 0 1086 160 6 N1END[1]
port 206 nsew signal input
rlabel metal2 s 1398 0 1454 160 6 N1END[2]
port 207 nsew signal input
rlabel metal2 s 1766 0 1822 160 6 N1END[3]
port 208 nsew signal input
rlabel metal2 s 2134 44840 2190 45000 6 N2BEG[0]
port 209 nsew signal output
rlabel metal2 s 2502 44840 2558 45000 6 N2BEG[1]
port 210 nsew signal output
rlabel metal2 s 2870 44840 2926 45000 6 N2BEG[2]
port 211 nsew signal output
rlabel metal2 s 3238 44840 3294 45000 6 N2BEG[3]
port 212 nsew signal output
rlabel metal2 s 3606 44840 3662 45000 6 N2BEG[4]
port 213 nsew signal output
rlabel metal2 s 3974 44840 4030 45000 6 N2BEG[5]
port 214 nsew signal output
rlabel metal2 s 4342 44840 4398 45000 6 N2BEG[6]
port 215 nsew signal output
rlabel metal2 s 4710 44840 4766 45000 6 N2BEG[7]
port 216 nsew signal output
rlabel metal2 s 5078 44840 5134 45000 6 N2BEGb[0]
port 217 nsew signal output
rlabel metal2 s 5446 44840 5502 45000 6 N2BEGb[1]
port 218 nsew signal output
rlabel metal2 s 5814 44840 5870 45000 6 N2BEGb[2]
port 219 nsew signal output
rlabel metal2 s 6182 44840 6238 45000 6 N2BEGb[3]
port 220 nsew signal output
rlabel metal2 s 6550 44840 6606 45000 6 N2BEGb[4]
port 221 nsew signal output
rlabel metal2 s 6918 44840 6974 45000 6 N2BEGb[5]
port 222 nsew signal output
rlabel metal2 s 7286 44840 7342 45000 6 N2BEGb[6]
port 223 nsew signal output
rlabel metal2 s 7654 44840 7710 45000 6 N2BEGb[7]
port 224 nsew signal output
rlabel metal2 s 5078 0 5134 160 6 N2END[0]
port 225 nsew signal input
rlabel metal2 s 5446 0 5502 160 6 N2END[1]
port 226 nsew signal input
rlabel metal2 s 5814 0 5870 160 6 N2END[2]
port 227 nsew signal input
rlabel metal2 s 6182 0 6238 160 6 N2END[3]
port 228 nsew signal input
rlabel metal2 s 6550 0 6606 160 6 N2END[4]
port 229 nsew signal input
rlabel metal2 s 6918 0 6974 160 6 N2END[5]
port 230 nsew signal input
rlabel metal2 s 7286 0 7342 160 6 N2END[6]
port 231 nsew signal input
rlabel metal2 s 7654 0 7710 160 6 N2END[7]
port 232 nsew signal input
rlabel metal2 s 2134 0 2190 160 6 N2MID[0]
port 233 nsew signal input
rlabel metal2 s 2502 0 2558 160 6 N2MID[1]
port 234 nsew signal input
rlabel metal2 s 2870 0 2926 160 6 N2MID[2]
port 235 nsew signal input
rlabel metal2 s 3238 0 3294 160 6 N2MID[3]
port 236 nsew signal input
rlabel metal2 s 3606 0 3662 160 6 N2MID[4]
port 237 nsew signal input
rlabel metal2 s 3974 0 4030 160 6 N2MID[5]
port 238 nsew signal input
rlabel metal2 s 4342 0 4398 160 6 N2MID[6]
port 239 nsew signal input
rlabel metal2 s 4710 0 4766 160 6 N2MID[7]
port 240 nsew signal input
rlabel metal2 s 8022 44840 8078 45000 6 N4BEG[0]
port 241 nsew signal output
rlabel metal2 s 11702 44840 11758 45000 6 N4BEG[10]
port 242 nsew signal output
rlabel metal2 s 12070 44840 12126 45000 6 N4BEG[11]
port 243 nsew signal output
rlabel metal2 s 12438 44840 12494 45000 6 N4BEG[12]
port 244 nsew signal output
rlabel metal2 s 12806 44840 12862 45000 6 N4BEG[13]
port 245 nsew signal output
rlabel metal2 s 13174 44840 13230 45000 6 N4BEG[14]
port 246 nsew signal output
rlabel metal2 s 13542 44840 13598 45000 6 N4BEG[15]
port 247 nsew signal output
rlabel metal2 s 8390 44840 8446 45000 6 N4BEG[1]
port 248 nsew signal output
rlabel metal2 s 8758 44840 8814 45000 6 N4BEG[2]
port 249 nsew signal output
rlabel metal2 s 9126 44840 9182 45000 6 N4BEG[3]
port 250 nsew signal output
rlabel metal2 s 9494 44840 9550 45000 6 N4BEG[4]
port 251 nsew signal output
rlabel metal2 s 9862 44840 9918 45000 6 N4BEG[5]
port 252 nsew signal output
rlabel metal2 s 10230 44840 10286 45000 6 N4BEG[6]
port 253 nsew signal output
rlabel metal2 s 10598 44840 10654 45000 6 N4BEG[7]
port 254 nsew signal output
rlabel metal2 s 10966 44840 11022 45000 6 N4BEG[8]
port 255 nsew signal output
rlabel metal2 s 11334 44840 11390 45000 6 N4BEG[9]
port 256 nsew signal output
rlabel metal2 s 8022 0 8078 160 6 N4END[0]
port 257 nsew signal input
rlabel metal2 s 11702 0 11758 160 6 N4END[10]
port 258 nsew signal input
rlabel metal2 s 12070 0 12126 160 6 N4END[11]
port 259 nsew signal input
rlabel metal2 s 12438 0 12494 160 6 N4END[12]
port 260 nsew signal input
rlabel metal2 s 12806 0 12862 160 6 N4END[13]
port 261 nsew signal input
rlabel metal2 s 13174 0 13230 160 6 N4END[14]
port 262 nsew signal input
rlabel metal2 s 13542 0 13598 160 6 N4END[15]
port 263 nsew signal input
rlabel metal2 s 8390 0 8446 160 6 N4END[1]
port 264 nsew signal input
rlabel metal2 s 8758 0 8814 160 6 N4END[2]
port 265 nsew signal input
rlabel metal2 s 9126 0 9182 160 6 N4END[3]
port 266 nsew signal input
rlabel metal2 s 9494 0 9550 160 6 N4END[4]
port 267 nsew signal input
rlabel metal2 s 9862 0 9918 160 6 N4END[5]
port 268 nsew signal input
rlabel metal2 s 10230 0 10286 160 6 N4END[6]
port 269 nsew signal input
rlabel metal2 s 10598 0 10654 160 6 N4END[7]
port 270 nsew signal input
rlabel metal2 s 10966 0 11022 160 6 N4END[8]
port 271 nsew signal input
rlabel metal2 s 11334 0 11390 160 6 N4END[9]
port 272 nsew signal input
rlabel metal2 s 13910 44840 13966 45000 6 NN4BEG[0]
port 273 nsew signal output
rlabel metal2 s 17590 44840 17646 45000 6 NN4BEG[10]
port 274 nsew signal output
rlabel metal2 s 17958 44840 18014 45000 6 NN4BEG[11]
port 275 nsew signal output
rlabel metal2 s 18326 44840 18382 45000 6 NN4BEG[12]
port 276 nsew signal output
rlabel metal2 s 18694 44840 18750 45000 6 NN4BEG[13]
port 277 nsew signal output
rlabel metal2 s 19062 44840 19118 45000 6 NN4BEG[14]
port 278 nsew signal output
rlabel metal2 s 19430 44840 19486 45000 6 NN4BEG[15]
port 279 nsew signal output
rlabel metal2 s 14278 44840 14334 45000 6 NN4BEG[1]
port 280 nsew signal output
rlabel metal2 s 14646 44840 14702 45000 6 NN4BEG[2]
port 281 nsew signal output
rlabel metal2 s 15014 44840 15070 45000 6 NN4BEG[3]
port 282 nsew signal output
rlabel metal2 s 15382 44840 15438 45000 6 NN4BEG[4]
port 283 nsew signal output
rlabel metal2 s 15750 44840 15806 45000 6 NN4BEG[5]
port 284 nsew signal output
rlabel metal2 s 16118 44840 16174 45000 6 NN4BEG[6]
port 285 nsew signal output
rlabel metal2 s 16486 44840 16542 45000 6 NN4BEG[7]
port 286 nsew signal output
rlabel metal2 s 16854 44840 16910 45000 6 NN4BEG[8]
port 287 nsew signal output
rlabel metal2 s 17222 44840 17278 45000 6 NN4BEG[9]
port 288 nsew signal output
rlabel metal2 s 13910 0 13966 160 6 NN4END[0]
port 289 nsew signal input
rlabel metal2 s 17590 0 17646 160 6 NN4END[10]
port 290 nsew signal input
rlabel metal2 s 17958 0 18014 160 6 NN4END[11]
port 291 nsew signal input
rlabel metal2 s 18326 0 18382 160 6 NN4END[12]
port 292 nsew signal input
rlabel metal2 s 18694 0 18750 160 6 NN4END[13]
port 293 nsew signal input
rlabel metal2 s 19062 0 19118 160 6 NN4END[14]
port 294 nsew signal input
rlabel metal2 s 19430 0 19486 160 6 NN4END[15]
port 295 nsew signal input
rlabel metal2 s 14278 0 14334 160 6 NN4END[1]
port 296 nsew signal input
rlabel metal2 s 14646 0 14702 160 6 NN4END[2]
port 297 nsew signal input
rlabel metal2 s 15014 0 15070 160 6 NN4END[3]
port 298 nsew signal input
rlabel metal2 s 15382 0 15438 160 6 NN4END[4]
port 299 nsew signal input
rlabel metal2 s 15750 0 15806 160 6 NN4END[5]
port 300 nsew signal input
rlabel metal2 s 16118 0 16174 160 6 NN4END[6]
port 301 nsew signal input
rlabel metal2 s 16486 0 16542 160 6 NN4END[7]
port 302 nsew signal input
rlabel metal2 s 16854 0 16910 160 6 NN4END[8]
port 303 nsew signal input
rlabel metal2 s 17222 0 17278 160 6 NN4END[9]
port 304 nsew signal input
rlabel metal2 s 19798 0 19854 160 6 S1BEG[0]
port 305 nsew signal output
rlabel metal2 s 20166 0 20222 160 6 S1BEG[1]
port 306 nsew signal output
rlabel metal2 s 20534 0 20590 160 6 S1BEG[2]
port 307 nsew signal output
rlabel metal2 s 20902 0 20958 160 6 S1BEG[3]
port 308 nsew signal output
rlabel metal2 s 19798 44840 19854 45000 6 S1END[0]
port 309 nsew signal input
rlabel metal2 s 20166 44840 20222 45000 6 S1END[1]
port 310 nsew signal input
rlabel metal2 s 20534 44840 20590 45000 6 S1END[2]
port 311 nsew signal input
rlabel metal2 s 20902 44840 20958 45000 6 S1END[3]
port 312 nsew signal input
rlabel metal2 s 24214 0 24270 160 6 S2BEG[0]
port 313 nsew signal output
rlabel metal2 s 24582 0 24638 160 6 S2BEG[1]
port 314 nsew signal output
rlabel metal2 s 24950 0 25006 160 6 S2BEG[2]
port 315 nsew signal output
rlabel metal2 s 25318 0 25374 160 6 S2BEG[3]
port 316 nsew signal output
rlabel metal2 s 25686 0 25742 160 6 S2BEG[4]
port 317 nsew signal output
rlabel metal2 s 26054 0 26110 160 6 S2BEG[5]
port 318 nsew signal output
rlabel metal2 s 26422 0 26478 160 6 S2BEG[6]
port 319 nsew signal output
rlabel metal2 s 26790 0 26846 160 6 S2BEG[7]
port 320 nsew signal output
rlabel metal2 s 21270 0 21326 160 6 S2BEGb[0]
port 321 nsew signal output
rlabel metal2 s 21638 0 21694 160 6 S2BEGb[1]
port 322 nsew signal output
rlabel metal2 s 22006 0 22062 160 6 S2BEGb[2]
port 323 nsew signal output
rlabel metal2 s 22374 0 22430 160 6 S2BEGb[3]
port 324 nsew signal output
rlabel metal2 s 22742 0 22798 160 6 S2BEGb[4]
port 325 nsew signal output
rlabel metal2 s 23110 0 23166 160 6 S2BEGb[5]
port 326 nsew signal output
rlabel metal2 s 23478 0 23534 160 6 S2BEGb[6]
port 327 nsew signal output
rlabel metal2 s 23846 0 23902 160 6 S2BEGb[7]
port 328 nsew signal output
rlabel metal2 s 21270 44840 21326 45000 6 S2END[0]
port 329 nsew signal input
rlabel metal2 s 21638 44840 21694 45000 6 S2END[1]
port 330 nsew signal input
rlabel metal2 s 22006 44840 22062 45000 6 S2END[2]
port 331 nsew signal input
rlabel metal2 s 22374 44840 22430 45000 6 S2END[3]
port 332 nsew signal input
rlabel metal2 s 22742 44840 22798 45000 6 S2END[4]
port 333 nsew signal input
rlabel metal2 s 23110 44840 23166 45000 6 S2END[5]
port 334 nsew signal input
rlabel metal2 s 23478 44840 23534 45000 6 S2END[6]
port 335 nsew signal input
rlabel metal2 s 23846 44840 23902 45000 6 S2END[7]
port 336 nsew signal input
rlabel metal2 s 24214 44840 24270 45000 6 S2MID[0]
port 337 nsew signal input
rlabel metal2 s 24582 44840 24638 45000 6 S2MID[1]
port 338 nsew signal input
rlabel metal2 s 24950 44840 25006 45000 6 S2MID[2]
port 339 nsew signal input
rlabel metal2 s 25318 44840 25374 45000 6 S2MID[3]
port 340 nsew signal input
rlabel metal2 s 25686 44840 25742 45000 6 S2MID[4]
port 341 nsew signal input
rlabel metal2 s 26054 44840 26110 45000 6 S2MID[5]
port 342 nsew signal input
rlabel metal2 s 26422 44840 26478 45000 6 S2MID[6]
port 343 nsew signal input
rlabel metal2 s 26790 44840 26846 45000 6 S2MID[7]
port 344 nsew signal input
rlabel metal2 s 27158 0 27214 160 6 S4BEG[0]
port 345 nsew signal output
rlabel metal2 s 30838 0 30894 160 6 S4BEG[10]
port 346 nsew signal output
rlabel metal2 s 31206 0 31262 160 6 S4BEG[11]
port 347 nsew signal output
rlabel metal2 s 31574 0 31630 160 6 S4BEG[12]
port 348 nsew signal output
rlabel metal2 s 31942 0 31998 160 6 S4BEG[13]
port 349 nsew signal output
rlabel metal2 s 32310 0 32366 160 6 S4BEG[14]
port 350 nsew signal output
rlabel metal2 s 32678 0 32734 160 6 S4BEG[15]
port 351 nsew signal output
rlabel metal2 s 27526 0 27582 160 6 S4BEG[1]
port 352 nsew signal output
rlabel metal2 s 27894 0 27950 160 6 S4BEG[2]
port 353 nsew signal output
rlabel metal2 s 28262 0 28318 160 6 S4BEG[3]
port 354 nsew signal output
rlabel metal2 s 28630 0 28686 160 6 S4BEG[4]
port 355 nsew signal output
rlabel metal2 s 28998 0 29054 160 6 S4BEG[5]
port 356 nsew signal output
rlabel metal2 s 29366 0 29422 160 6 S4BEG[6]
port 357 nsew signal output
rlabel metal2 s 29734 0 29790 160 6 S4BEG[7]
port 358 nsew signal output
rlabel metal2 s 30102 0 30158 160 6 S4BEG[8]
port 359 nsew signal output
rlabel metal2 s 30470 0 30526 160 6 S4BEG[9]
port 360 nsew signal output
rlabel metal2 s 27158 44840 27214 45000 6 S4END[0]
port 361 nsew signal input
rlabel metal2 s 30838 44840 30894 45000 6 S4END[10]
port 362 nsew signal input
rlabel metal2 s 31206 44840 31262 45000 6 S4END[11]
port 363 nsew signal input
rlabel metal2 s 31574 44840 31630 45000 6 S4END[12]
port 364 nsew signal input
rlabel metal2 s 31942 44840 31998 45000 6 S4END[13]
port 365 nsew signal input
rlabel metal2 s 32310 44840 32366 45000 6 S4END[14]
port 366 nsew signal input
rlabel metal2 s 32678 44840 32734 45000 6 S4END[15]
port 367 nsew signal input
rlabel metal2 s 27526 44840 27582 45000 6 S4END[1]
port 368 nsew signal input
rlabel metal2 s 27894 44840 27950 45000 6 S4END[2]
port 369 nsew signal input
rlabel metal2 s 28262 44840 28318 45000 6 S4END[3]
port 370 nsew signal input
rlabel metal2 s 28630 44840 28686 45000 6 S4END[4]
port 371 nsew signal input
rlabel metal2 s 28998 44840 29054 45000 6 S4END[5]
port 372 nsew signal input
rlabel metal2 s 29366 44840 29422 45000 6 S4END[6]
port 373 nsew signal input
rlabel metal2 s 29734 44840 29790 45000 6 S4END[7]
port 374 nsew signal input
rlabel metal2 s 30102 44840 30158 45000 6 S4END[8]
port 375 nsew signal input
rlabel metal2 s 30470 44840 30526 45000 6 S4END[9]
port 376 nsew signal input
rlabel metal2 s 33046 0 33102 160 6 SS4BEG[0]
port 377 nsew signal output
rlabel metal2 s 36726 0 36782 160 6 SS4BEG[10]
port 378 nsew signal output
rlabel metal2 s 37094 0 37150 160 6 SS4BEG[11]
port 379 nsew signal output
rlabel metal2 s 37462 0 37518 160 6 SS4BEG[12]
port 380 nsew signal output
rlabel metal2 s 37830 0 37886 160 6 SS4BEG[13]
port 381 nsew signal output
rlabel metal2 s 38198 0 38254 160 6 SS4BEG[14]
port 382 nsew signal output
rlabel metal2 s 38566 0 38622 160 6 SS4BEG[15]
port 383 nsew signal output
rlabel metal2 s 33414 0 33470 160 6 SS4BEG[1]
port 384 nsew signal output
rlabel metal2 s 33782 0 33838 160 6 SS4BEG[2]
port 385 nsew signal output
rlabel metal2 s 34150 0 34206 160 6 SS4BEG[3]
port 386 nsew signal output
rlabel metal2 s 34518 0 34574 160 6 SS4BEG[4]
port 387 nsew signal output
rlabel metal2 s 34886 0 34942 160 6 SS4BEG[5]
port 388 nsew signal output
rlabel metal2 s 35254 0 35310 160 6 SS4BEG[6]
port 389 nsew signal output
rlabel metal2 s 35622 0 35678 160 6 SS4BEG[7]
port 390 nsew signal output
rlabel metal2 s 35990 0 36046 160 6 SS4BEG[8]
port 391 nsew signal output
rlabel metal2 s 36358 0 36414 160 6 SS4BEG[9]
port 392 nsew signal output
rlabel metal2 s 33046 44840 33102 45000 6 SS4END[0]
port 393 nsew signal input
rlabel metal2 s 36726 44840 36782 45000 6 SS4END[10]
port 394 nsew signal input
rlabel metal2 s 37094 44840 37150 45000 6 SS4END[11]
port 395 nsew signal input
rlabel metal2 s 37462 44840 37518 45000 6 SS4END[12]
port 396 nsew signal input
rlabel metal2 s 37830 44840 37886 45000 6 SS4END[13]
port 397 nsew signal input
rlabel metal2 s 38198 44840 38254 45000 6 SS4END[14]
port 398 nsew signal input
rlabel metal2 s 38566 44840 38622 45000 6 SS4END[15]
port 399 nsew signal input
rlabel metal2 s 33414 44840 33470 45000 6 SS4END[1]
port 400 nsew signal input
rlabel metal2 s 33782 44840 33838 45000 6 SS4END[2]
port 401 nsew signal input
rlabel metal2 s 34150 44840 34206 45000 6 SS4END[3]
port 402 nsew signal input
rlabel metal2 s 34518 44840 34574 45000 6 SS4END[4]
port 403 nsew signal input
rlabel metal2 s 34886 44840 34942 45000 6 SS4END[5]
port 404 nsew signal input
rlabel metal2 s 35254 44840 35310 45000 6 SS4END[6]
port 405 nsew signal input
rlabel metal2 s 35622 44840 35678 45000 6 SS4END[7]
port 406 nsew signal input
rlabel metal2 s 35990 44840 36046 45000 6 SS4END[8]
port 407 nsew signal input
rlabel metal2 s 36358 44840 36414 45000 6 SS4END[9]
port 408 nsew signal input
rlabel metal2 s 38934 0 38990 160 6 UserCLK
port 409 nsew signal input
rlabel metal2 s 38934 44840 38990 45000 6 UserCLKo
port 410 nsew signal output
rlabel metal4 s 19568 1040 19888 43568 6 VGND
port 411 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 43568 6 VPWR
port 412 nsew power bidirectional
rlabel metal4 s 34928 1040 35248 43568 6 VPWR
port 412 nsew power bidirectional
rlabel metal3 s 0 5176 160 5296 6 W1BEG[0]
port 413 nsew signal output
rlabel metal3 s 0 5448 160 5568 6 W1BEG[1]
port 414 nsew signal output
rlabel metal3 s 0 5720 160 5840 6 W1BEG[2]
port 415 nsew signal output
rlabel metal3 s 0 5992 160 6112 6 W1BEG[3]
port 416 nsew signal output
rlabel metal3 s 46840 5176 47000 5296 6 W1END[0]
port 417 nsew signal input
rlabel metal3 s 46840 5448 47000 5568 6 W1END[1]
port 418 nsew signal input
rlabel metal3 s 46840 5720 47000 5840 6 W1END[2]
port 419 nsew signal input
rlabel metal3 s 46840 5992 47000 6112 6 W1END[3]
port 420 nsew signal input
rlabel metal3 s 0 6264 160 6384 6 W2BEG[0]
port 421 nsew signal output
rlabel metal3 s 0 6536 160 6656 6 W2BEG[1]
port 422 nsew signal output
rlabel metal3 s 0 6808 160 6928 6 W2BEG[2]
port 423 nsew signal output
rlabel metal3 s 0 7080 160 7200 6 W2BEG[3]
port 424 nsew signal output
rlabel metal3 s 0 7352 160 7472 6 W2BEG[4]
port 425 nsew signal output
rlabel metal3 s 0 7624 160 7744 6 W2BEG[5]
port 426 nsew signal output
rlabel metal3 s 0 7896 160 8016 6 W2BEG[6]
port 427 nsew signal output
rlabel metal3 s 0 8168 160 8288 6 W2BEG[7]
port 428 nsew signal output
rlabel metal3 s 0 8440 160 8560 6 W2BEGb[0]
port 429 nsew signal output
rlabel metal3 s 0 8712 160 8832 6 W2BEGb[1]
port 430 nsew signal output
rlabel metal3 s 0 8984 160 9104 6 W2BEGb[2]
port 431 nsew signal output
rlabel metal3 s 0 9256 160 9376 6 W2BEGb[3]
port 432 nsew signal output
rlabel metal3 s 0 9528 160 9648 6 W2BEGb[4]
port 433 nsew signal output
rlabel metal3 s 0 9800 160 9920 6 W2BEGb[5]
port 434 nsew signal output
rlabel metal3 s 0 10072 160 10192 6 W2BEGb[6]
port 435 nsew signal output
rlabel metal3 s 0 10344 160 10464 6 W2BEGb[7]
port 436 nsew signal output
rlabel metal3 s 46840 8440 47000 8560 6 W2END[0]
port 437 nsew signal input
rlabel metal3 s 46840 8712 47000 8832 6 W2END[1]
port 438 nsew signal input
rlabel metal3 s 46840 8984 47000 9104 6 W2END[2]
port 439 nsew signal input
rlabel metal3 s 46840 9256 47000 9376 6 W2END[3]
port 440 nsew signal input
rlabel metal3 s 46840 9528 47000 9648 6 W2END[4]
port 441 nsew signal input
rlabel metal3 s 46840 9800 47000 9920 6 W2END[5]
port 442 nsew signal input
rlabel metal3 s 46840 10072 47000 10192 6 W2END[6]
port 443 nsew signal input
rlabel metal3 s 46840 10344 47000 10464 6 W2END[7]
port 444 nsew signal input
rlabel metal3 s 46840 6264 47000 6384 6 W2MID[0]
port 445 nsew signal input
rlabel metal3 s 46840 6536 47000 6656 6 W2MID[1]
port 446 nsew signal input
rlabel metal3 s 46840 6808 47000 6928 6 W2MID[2]
port 447 nsew signal input
rlabel metal3 s 46840 7080 47000 7200 6 W2MID[3]
port 448 nsew signal input
rlabel metal3 s 46840 7352 47000 7472 6 W2MID[4]
port 449 nsew signal input
rlabel metal3 s 46840 7624 47000 7744 6 W2MID[5]
port 450 nsew signal input
rlabel metal3 s 46840 7896 47000 8016 6 W2MID[6]
port 451 nsew signal input
rlabel metal3 s 46840 8168 47000 8288 6 W2MID[7]
port 452 nsew signal input
rlabel metal3 s 0 14968 160 15088 6 W6BEG[0]
port 453 nsew signal output
rlabel metal3 s 0 17688 160 17808 6 W6BEG[10]
port 454 nsew signal output
rlabel metal3 s 0 17960 160 18080 6 W6BEG[11]
port 455 nsew signal output
rlabel metal3 s 0 15240 160 15360 6 W6BEG[1]
port 456 nsew signal output
rlabel metal3 s 0 15512 160 15632 6 W6BEG[2]
port 457 nsew signal output
rlabel metal3 s 0 15784 160 15904 6 W6BEG[3]
port 458 nsew signal output
rlabel metal3 s 0 16056 160 16176 6 W6BEG[4]
port 459 nsew signal output
rlabel metal3 s 0 16328 160 16448 6 W6BEG[5]
port 460 nsew signal output
rlabel metal3 s 0 16600 160 16720 6 W6BEG[6]
port 461 nsew signal output
rlabel metal3 s 0 16872 160 16992 6 W6BEG[7]
port 462 nsew signal output
rlabel metal3 s 0 17144 160 17264 6 W6BEG[8]
port 463 nsew signal output
rlabel metal3 s 0 17416 160 17536 6 W6BEG[9]
port 464 nsew signal output
rlabel metal3 s 46840 14968 47000 15088 6 W6END[0]
port 465 nsew signal input
rlabel metal3 s 46840 17688 47000 17808 6 W6END[10]
port 466 nsew signal input
rlabel metal3 s 46840 17960 47000 18080 6 W6END[11]
port 467 nsew signal input
rlabel metal3 s 46840 15240 47000 15360 6 W6END[1]
port 468 nsew signal input
rlabel metal3 s 46840 15512 47000 15632 6 W6END[2]
port 469 nsew signal input
rlabel metal3 s 46840 15784 47000 15904 6 W6END[3]
port 470 nsew signal input
rlabel metal3 s 46840 16056 47000 16176 6 W6END[4]
port 471 nsew signal input
rlabel metal3 s 46840 16328 47000 16448 6 W6END[5]
port 472 nsew signal input
rlabel metal3 s 46840 16600 47000 16720 6 W6END[6]
port 473 nsew signal input
rlabel metal3 s 46840 16872 47000 16992 6 W6END[7]
port 474 nsew signal input
rlabel metal3 s 46840 17144 47000 17264 6 W6END[8]
port 475 nsew signal input
rlabel metal3 s 46840 17416 47000 17536 6 W6END[9]
port 476 nsew signal input
rlabel metal3 s 0 10616 160 10736 6 WW4BEG[0]
port 477 nsew signal output
rlabel metal3 s 0 13336 160 13456 6 WW4BEG[10]
port 478 nsew signal output
rlabel metal3 s 0 13608 160 13728 6 WW4BEG[11]
port 479 nsew signal output
rlabel metal3 s 0 13880 160 14000 6 WW4BEG[12]
port 480 nsew signal output
rlabel metal3 s 0 14152 160 14272 6 WW4BEG[13]
port 481 nsew signal output
rlabel metal3 s 0 14424 160 14544 6 WW4BEG[14]
port 482 nsew signal output
rlabel metal3 s 0 14696 160 14816 6 WW4BEG[15]
port 483 nsew signal output
rlabel metal3 s 0 10888 160 11008 6 WW4BEG[1]
port 484 nsew signal output
rlabel metal3 s 0 11160 160 11280 6 WW4BEG[2]
port 485 nsew signal output
rlabel metal3 s 0 11432 160 11552 6 WW4BEG[3]
port 486 nsew signal output
rlabel metal3 s 0 11704 160 11824 6 WW4BEG[4]
port 487 nsew signal output
rlabel metal3 s 0 11976 160 12096 6 WW4BEG[5]
port 488 nsew signal output
rlabel metal3 s 0 12248 160 12368 6 WW4BEG[6]
port 489 nsew signal output
rlabel metal3 s 0 12520 160 12640 6 WW4BEG[7]
port 490 nsew signal output
rlabel metal3 s 0 12792 160 12912 6 WW4BEG[8]
port 491 nsew signal output
rlabel metal3 s 0 13064 160 13184 6 WW4BEG[9]
port 492 nsew signal output
rlabel metal3 s 46840 10616 47000 10736 6 WW4END[0]
port 493 nsew signal input
rlabel metal3 s 46840 13336 47000 13456 6 WW4END[10]
port 494 nsew signal input
rlabel metal3 s 46840 13608 47000 13728 6 WW4END[11]
port 495 nsew signal input
rlabel metal3 s 46840 13880 47000 14000 6 WW4END[12]
port 496 nsew signal input
rlabel metal3 s 46840 14152 47000 14272 6 WW4END[13]
port 497 nsew signal input
rlabel metal3 s 46840 14424 47000 14544 6 WW4END[14]
port 498 nsew signal input
rlabel metal3 s 46840 14696 47000 14816 6 WW4END[15]
port 499 nsew signal input
rlabel metal3 s 46840 10888 47000 11008 6 WW4END[1]
port 500 nsew signal input
rlabel metal3 s 46840 11160 47000 11280 6 WW4END[2]
port 501 nsew signal input
rlabel metal3 s 46840 11432 47000 11552 6 WW4END[3]
port 502 nsew signal input
rlabel metal3 s 46840 11704 47000 11824 6 WW4END[4]
port 503 nsew signal input
rlabel metal3 s 46840 11976 47000 12096 6 WW4END[5]
port 504 nsew signal input
rlabel metal3 s 46840 12248 47000 12368 6 WW4END[6]
port 505 nsew signal input
rlabel metal3 s 46840 12520 47000 12640 6 WW4END[7]
port 506 nsew signal input
rlabel metal3 s 46840 12792 47000 12912 6 WW4END[8]
port 507 nsew signal input
rlabel metal3 s 46840 13064 47000 13184 6 WW4END[9]
port 508 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 47000 45000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7634980
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/RegFile/runs/24_12_05_10_24/results/signoff/RegFile.magic.gds
string GDS_START 275338
<< end >>

