magic
tech sky130A
magscale 1 2
timestamp 1733268178
<< viali >>
rect 2053 8585 2087 8619
rect 2789 8585 2823 8619
rect 3157 8585 3191 8619
rect 4261 8585 4295 8619
rect 4813 8585 4847 8619
rect 5365 8585 5399 8619
rect 5733 8585 5767 8619
rect 6653 8585 6687 8619
rect 7389 8585 7423 8619
rect 7757 8585 7791 8619
rect 8309 8585 8343 8619
rect 8677 8585 8711 8619
rect 9229 8585 9263 8619
rect 9597 8585 9631 8619
rect 12081 8585 12115 8619
rect 12357 8585 12391 8619
rect 13093 8585 13127 8619
rect 13921 8585 13955 8619
rect 14381 8585 14415 8619
rect 15209 8585 15243 8619
rect 15761 8585 15795 8619
rect 15853 8585 15887 8619
rect 16129 8585 16163 8619
rect 16681 8585 16715 8619
rect 16957 8585 16991 8619
rect 17233 8585 17267 8619
rect 17509 8585 17543 8619
rect 19073 8585 19107 8619
rect 19993 8585 20027 8619
rect 20361 8585 20395 8619
rect 20729 8585 20763 8619
rect 21281 8585 21315 8619
rect 22385 8585 22419 8619
rect 22937 8585 22971 8619
rect 23489 8585 23523 8619
rect 3985 8517 4019 8551
rect 5089 8517 5123 8551
rect 8033 8517 8067 8551
rect 1961 8449 1995 8483
rect 2513 8449 2547 8483
rect 3065 8449 3099 8483
rect 4629 8449 4663 8483
rect 5641 8449 5675 8483
rect 6561 8449 6595 8483
rect 7205 8449 7239 8483
rect 7573 8449 7607 8483
rect 8493 8449 8527 8483
rect 9045 8449 9079 8483
rect 9413 8449 9447 8483
rect 10057 8449 10091 8483
rect 10241 8449 10275 8483
rect 10701 8449 10735 8483
rect 11345 8449 11379 8483
rect 11713 8449 11747 8483
rect 11989 8449 12023 8483
rect 12265 8449 12299 8483
rect 12541 8453 12575 8487
rect 12633 8449 12667 8483
rect 12909 8449 12943 8483
rect 13369 8449 13403 8483
rect 13645 8449 13679 8483
rect 13737 8449 13771 8483
rect 14197 8449 14231 8483
rect 14657 8449 14691 8483
rect 14933 8449 14967 8483
rect 15025 8449 15059 8483
rect 15485 8449 15519 8483
rect 15577 8449 15611 8483
rect 16037 8449 16071 8483
rect 16313 8449 16347 8483
rect 16865 8449 16899 8483
rect 17141 8449 17175 8483
rect 17417 8449 17451 8483
rect 17693 8449 17727 8483
rect 17785 8449 17819 8483
rect 18061 8449 18095 8483
rect 18521 8449 18555 8483
rect 18797 8449 18831 8483
rect 18889 8449 18923 8483
rect 19441 8449 19475 8483
rect 19717 8449 19751 8483
rect 19809 8449 19843 8483
rect 20177 8449 20211 8483
rect 20637 8449 20671 8483
rect 21189 8449 21223 8483
rect 21833 8449 21867 8483
rect 22293 8449 22327 8483
rect 22845 8449 22879 8483
rect 23397 8449 23431 8483
rect 10425 8313 10459 8347
rect 10885 8313 10919 8347
rect 11529 8313 11563 8347
rect 13185 8313 13219 8347
rect 13461 8313 13495 8347
rect 14473 8313 14507 8347
rect 15301 8313 15335 8347
rect 17969 8313 18003 8347
rect 18245 8313 18279 8347
rect 18337 8313 18371 8347
rect 22017 8313 22051 8347
rect 9873 8245 9907 8279
rect 11161 8245 11195 8279
rect 11805 8245 11839 8279
rect 12817 8245 12851 8279
rect 14749 8245 14783 8279
rect 18613 8245 18647 8279
rect 19257 8245 19291 8279
rect 19533 8245 19567 8279
rect 1685 8041 1719 8075
rect 2421 8041 2455 8075
rect 2789 8041 2823 8075
rect 3341 8041 3375 8075
rect 4169 8041 4203 8075
rect 4997 8041 5031 8075
rect 6101 8041 6135 8075
rect 6653 8041 6687 8075
rect 7205 8041 7239 8075
rect 7757 8041 7791 8075
rect 8309 8041 8343 8075
rect 11069 8041 11103 8075
rect 11621 8041 11655 8075
rect 13001 8041 13035 8075
rect 14933 8041 14967 8075
rect 15209 8041 15243 8075
rect 15853 8041 15887 8075
rect 16405 8041 16439 8075
rect 16957 8041 16991 8075
rect 17509 8041 17543 8075
rect 17969 8041 18003 8075
rect 21097 8041 21131 8075
rect 22569 8041 22603 8075
rect 23121 8041 23155 8075
rect 23949 8041 23983 8075
rect 5733 7973 5767 8007
rect 9413 7973 9447 8007
rect 9873 7973 9907 8007
rect 11345 7973 11379 8007
rect 12449 7973 12483 8007
rect 13277 7973 13311 8007
rect 15577 7973 15611 8007
rect 16129 7973 16163 8007
rect 17233 7973 17267 8007
rect 18245 7973 18279 8007
rect 18981 7973 19015 8007
rect 22201 7973 22235 8007
rect 1593 7837 1627 7871
rect 2145 7837 2179 7871
rect 2697 7837 2731 7871
rect 3249 7837 3283 7871
rect 4077 7837 4111 7871
rect 5549 7837 5583 7871
rect 7573 7837 7607 7871
rect 8217 7837 8251 7871
rect 9321 7837 9355 7871
rect 9597 7837 9631 7871
rect 9689 7853 9723 7887
rect 10149 7837 10183 7871
rect 10425 7837 10459 7871
rect 10701 7837 10735 7871
rect 10977 7837 11011 7871
rect 11253 7837 11287 7871
rect 11529 7837 11563 7871
rect 11805 7837 11839 7871
rect 12081 7837 12115 7871
rect 12633 7837 12667 7871
rect 13185 7837 13219 7871
rect 13461 7837 13495 7871
rect 15117 7837 15151 7871
rect 15393 7837 15427 7871
rect 15761 7837 15795 7871
rect 16037 7837 16071 7871
rect 16313 7837 16347 7871
rect 16589 7837 16623 7871
rect 16865 7837 16899 7871
rect 17141 7837 17175 7871
rect 17417 7837 17451 7871
rect 17693 7837 17727 7871
rect 17785 7837 17819 7871
rect 18429 7837 18463 7871
rect 18521 7837 18555 7871
rect 18797 7837 18831 7871
rect 19349 7837 19383 7871
rect 19625 7837 19659 7871
rect 19901 7837 19935 7871
rect 20913 7837 20947 7871
rect 21741 7837 21775 7871
rect 4905 7769 4939 7803
rect 6009 7769 6043 7803
rect 6561 7769 6595 7803
rect 7113 7769 7147 7803
rect 21373 7769 21407 7803
rect 21925 7769 21959 7803
rect 22477 7769 22511 7803
rect 23029 7769 23063 7803
rect 23857 7769 23891 7803
rect 9137 7701 9171 7735
rect 9965 7701 9999 7735
rect 10241 7701 10275 7735
rect 10517 7701 10551 7735
rect 10793 7701 10827 7735
rect 11897 7701 11931 7735
rect 16681 7701 16715 7735
rect 18705 7701 18739 7735
rect 19533 7701 19567 7735
rect 19809 7701 19843 7735
rect 20085 7701 20119 7735
rect 2053 7497 2087 7531
rect 2789 7497 2823 7531
rect 3525 7497 3559 7531
rect 4629 7497 4663 7531
rect 5457 7497 5491 7531
rect 5733 7497 5767 7531
rect 6009 7497 6043 7531
rect 6653 7497 6687 7531
rect 7481 7497 7515 7531
rect 7757 7497 7791 7531
rect 8033 7497 8067 7531
rect 8585 7497 8619 7531
rect 10241 7497 10275 7531
rect 22293 7497 22327 7531
rect 23949 7497 23983 7531
rect 1961 7429 1995 7463
rect 2513 7429 2547 7463
rect 22937 7429 22971 7463
rect 2973 7361 3007 7395
rect 3341 7361 3375 7395
rect 4445 7361 4479 7395
rect 5641 7361 5675 7395
rect 5917 7361 5951 7395
rect 6193 7361 6227 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 7205 7361 7239 7395
rect 7665 7361 7699 7395
rect 7941 7361 7975 7395
rect 8217 7361 8251 7395
rect 8769 7361 8803 7395
rect 10425 7361 10459 7395
rect 22017 7361 22051 7395
rect 22569 7361 22603 7395
rect 23121 7361 23155 7395
rect 23673 7361 23707 7395
rect 23397 7293 23431 7327
rect 3157 7157 3191 7191
rect 6377 7157 6411 7191
rect 23121 6953 23155 6987
rect 1961 6817 1995 6851
rect 23949 6817 23983 6851
rect 1685 6749 1719 6783
rect 23673 6749 23707 6783
rect 2237 6681 2271 6715
rect 23029 6681 23063 6715
rect 2329 6613 2363 6647
rect 1593 6409 1627 6443
rect 23765 6409 23799 6443
rect 24317 6409 24351 6443
rect 1501 6341 1535 6375
rect 24041 6341 24075 6375
rect 17509 6273 17543 6307
rect 23489 6273 23523 6307
rect 17325 6069 17359 6103
rect 16773 5865 16807 5899
rect 16957 5661 16991 5695
rect 9137 2057 9171 2091
rect 10241 2057 10275 2091
rect 10609 2057 10643 2091
rect 11713 2057 11747 2091
rect 12817 2057 12851 2091
rect 13093 2057 13127 2091
rect 13829 2057 13863 2091
rect 15117 2057 15151 2091
rect 16313 2057 16347 2091
rect 20361 2057 20395 2091
rect 22109 2057 22143 2091
rect 22385 2057 22419 2091
rect 23581 2057 23615 2091
rect 23857 2057 23891 2091
rect 24133 2057 24167 2091
rect 7757 1921 7791 1955
rect 8953 1921 8987 1955
rect 10057 1921 10091 1955
rect 10425 1921 10459 1955
rect 11529 1921 11563 1955
rect 12633 1921 12667 1955
rect 12909 1921 12943 1955
rect 13645 1921 13679 1955
rect 13921 1921 13955 1955
rect 14933 1921 14967 1955
rect 15393 1921 15427 1955
rect 16129 1921 16163 1955
rect 18613 1921 18647 1955
rect 20545 1921 20579 1955
rect 22293 1921 22327 1955
rect 22569 1921 22603 1955
rect 23489 1921 23523 1955
rect 23765 1921 23799 1955
rect 24041 1921 24075 1955
rect 24317 1921 24351 1955
rect 7941 1785 7975 1819
rect 14105 1785 14139 1819
rect 18797 1785 18831 1819
rect 15577 1717 15611 1751
rect 23305 1717 23339 1751
rect 7205 1513 7239 1547
rect 8401 1513 8435 1547
rect 9597 1513 9631 1547
rect 9873 1513 9907 1547
rect 10885 1513 10919 1547
rect 12357 1513 12391 1547
rect 13185 1513 13219 1547
rect 14473 1513 14507 1547
rect 15669 1513 15703 1547
rect 18153 1513 18187 1547
rect 20177 1513 20211 1547
rect 21833 1513 21867 1547
rect 22845 1513 22879 1547
rect 23765 1513 23799 1547
rect 13461 1445 13495 1479
rect 21373 1445 21407 1479
rect 22109 1445 22143 1479
rect 23489 1445 23523 1479
rect 1409 1309 1443 1343
rect 2237 1309 2271 1343
rect 3433 1309 3467 1343
rect 4813 1309 4847 1343
rect 6009 1309 6043 1343
rect 7389 1309 7423 1343
rect 7665 1309 7699 1343
rect 8585 1309 8619 1343
rect 9137 1309 9171 1343
rect 9781 1309 9815 1343
rect 10057 1309 10091 1343
rect 10333 1309 10367 1343
rect 10793 1309 10827 1343
rect 11069 1309 11103 1343
rect 11989 1309 12023 1343
rect 12265 1309 12299 1343
rect 12541 1309 12575 1343
rect 13369 1309 13403 1343
rect 13645 1309 13679 1343
rect 13921 1309 13955 1343
rect 14381 1309 14415 1343
rect 14657 1309 14691 1343
rect 15025 1309 15059 1343
rect 15577 1309 15611 1343
rect 15853 1309 15887 1343
rect 16681 1309 16715 1343
rect 17141 1309 17175 1343
rect 17969 1309 18003 1343
rect 18337 1309 18371 1343
rect 19441 1309 19475 1343
rect 20361 1309 20395 1343
rect 21557 1309 21591 1343
rect 22017 1309 22051 1343
rect 22293 1309 22327 1343
rect 22753 1309 22787 1343
rect 23029 1309 23063 1343
rect 23397 1309 23431 1343
rect 23673 1309 23707 1343
rect 23949 1309 23983 1343
rect 24225 1309 24259 1343
rect 1593 1173 1627 1207
rect 2421 1173 2455 1207
rect 3617 1173 3651 1207
rect 4629 1173 4663 1207
rect 5825 1173 5859 1207
rect 7481 1173 7515 1207
rect 8953 1173 8987 1207
rect 10149 1173 10183 1207
rect 10609 1173 10643 1207
rect 11805 1173 11839 1207
rect 12081 1173 12115 1207
rect 13737 1173 13771 1207
rect 14197 1173 14231 1207
rect 14841 1173 14875 1207
rect 15393 1173 15427 1207
rect 16865 1173 16899 1207
rect 16957 1173 16991 1207
rect 17785 1173 17819 1207
rect 19257 1173 19291 1207
rect 22569 1173 22603 1207
rect 23213 1173 23247 1207
rect 24041 1173 24075 1207
<< metal1 >>
rect 7834 9936 7840 9988
rect 7892 9976 7898 9988
rect 18598 9976 18604 9988
rect 7892 9948 18604 9976
rect 7892 9936 7898 9948
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 18506 9908 18512 9920
rect 6656 9880 18512 9908
rect 6656 9784 6684 9880
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 15010 9840 15016 9852
rect 7484 9812 15016 9840
rect 7484 9784 7512 9812
rect 15010 9800 15016 9812
rect 15068 9800 15074 9852
rect 6638 9732 6644 9784
rect 6696 9732 6702 9784
rect 7466 9732 7472 9784
rect 7524 9732 7530 9784
rect 10594 9732 10600 9784
rect 10652 9772 10658 9784
rect 14090 9772 14096 9784
rect 10652 9744 14096 9772
rect 10652 9732 10658 9744
rect 14090 9732 14096 9744
rect 14148 9732 14154 9784
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 15194 9704 15200 9716
rect 3752 9676 15200 9704
rect 3752 9664 3758 9676
rect 15194 9664 15200 9676
rect 15252 9664 15258 9716
rect 7558 9596 7564 9648
rect 7616 9636 7622 9648
rect 18230 9636 18236 9648
rect 7616 9608 18236 9636
rect 7616 9596 7622 9608
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 11606 9568 11612 9580
rect 2924 9540 11612 9568
rect 2924 9528 2930 9540
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 11698 9528 11704 9580
rect 11756 9568 11762 9580
rect 19978 9568 19984 9580
rect 11756 9540 19984 9568
rect 11756 9528 11762 9540
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 8938 9460 8944 9512
rect 8996 9500 9002 9512
rect 16298 9500 16304 9512
rect 8996 9472 16304 9500
rect 8996 9460 9002 9472
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 8386 9392 8392 9444
rect 8444 9432 8450 9444
rect 13538 9432 13544 9444
rect 8444 9404 13544 9432
rect 8444 9392 8450 9404
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 2498 9324 2504 9376
rect 2556 9364 2562 9376
rect 11422 9364 11428 9376
rect 2556 9336 11428 9364
rect 2556 9324 2562 9336
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 14182 9364 14188 9376
rect 11664 9336 14188 9364
rect 11664 9324 11670 9336
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 2774 9256 2780 9308
rect 2832 9296 2838 9308
rect 13906 9296 13912 9308
rect 2832 9268 13912 9296
rect 2832 9256 2838 9268
rect 13906 9256 13912 9268
rect 13964 9256 13970 9308
rect 2314 9188 2320 9240
rect 2372 9228 2378 9240
rect 2372 9200 3924 9228
rect 2372 9188 2378 9200
rect 1762 9120 1768 9172
rect 1820 9160 1826 9172
rect 3694 9160 3700 9172
rect 1820 9132 3700 9160
rect 1820 9120 1826 9132
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 3896 9160 3924 9200
rect 8018 9188 8024 9240
rect 8076 9228 8082 9240
rect 17494 9228 17500 9240
rect 8076 9200 17500 9228
rect 8076 9188 8082 9200
rect 17494 9188 17500 9200
rect 17552 9188 17558 9240
rect 12618 9160 12624 9172
rect 3896 9132 12624 9160
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 19702 9160 19708 9172
rect 18748 9132 19708 9160
rect 18748 9120 18754 9132
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 9398 9052 9404 9104
rect 9456 9092 9462 9104
rect 16666 9092 16672 9104
rect 9456 9064 16672 9092
rect 9456 9052 9462 9064
rect 16666 9052 16672 9064
rect 16724 9052 16730 9104
rect 21726 9052 21732 9104
rect 21784 9092 21790 9104
rect 22922 9092 22928 9104
rect 21784 9064 22928 9092
rect 21784 9052 21790 9064
rect 22922 9052 22928 9064
rect 22980 9052 22986 9104
rect 16942 9024 16948 9036
rect 9232 8996 16948 9024
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 8662 8888 8668 8900
rect 5592 8860 8668 8888
rect 5592 8848 5598 8860
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 9232 8832 9260 8996
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17218 8956 17224 8968
rect 9968 8928 17224 8956
rect 9968 8832 9996 8928
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 15838 8888 15844 8900
rect 11164 8860 15844 8888
rect 11164 8832 11192 8860
rect 15838 8848 15844 8860
rect 15896 8848 15902 8900
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 8386 8820 8392 8832
rect 3200 8792 8392 8820
rect 3200 8780 3206 8792
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 9214 8780 9220 8832
rect 9272 8780 9278 8832
rect 9950 8780 9956 8832
rect 10008 8780 10014 8832
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 12710 8780 12716 8832
rect 12768 8820 12774 8832
rect 14734 8820 14740 8832
rect 12768 8792 14740 8820
rect 12768 8780 12774 8792
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 1104 8730 25000 8752
rect 1104 8678 6884 8730
rect 6936 8678 6948 8730
rect 7000 8678 7012 8730
rect 7064 8678 7076 8730
rect 7128 8678 7140 8730
rect 7192 8678 12818 8730
rect 12870 8678 12882 8730
rect 12934 8678 12946 8730
rect 12998 8678 13010 8730
rect 13062 8678 13074 8730
rect 13126 8678 18752 8730
rect 18804 8678 18816 8730
rect 18868 8678 18880 8730
rect 18932 8678 18944 8730
rect 18996 8678 19008 8730
rect 19060 8678 24686 8730
rect 24738 8678 24750 8730
rect 24802 8678 24814 8730
rect 24866 8678 24878 8730
rect 24930 8678 24942 8730
rect 24994 8678 25000 8730
rect 1104 8656 25000 8678
rect 2038 8576 2044 8628
rect 2096 8576 2102 8628
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 2958 8616 2964 8628
rect 2823 8588 2964 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 3145 8619 3203 8625
rect 3145 8585 3157 8619
rect 3191 8585 3203 8619
rect 3145 8579 3203 8585
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4338 8616 4344 8628
rect 4295 8588 4344 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 658 8508 664 8560
rect 716 8548 722 8560
rect 3160 8548 3188 8579
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4801 8619 4859 8625
rect 4801 8585 4813 8619
rect 4847 8616 4859 8619
rect 5166 8616 5172 8628
rect 4847 8588 5172 8616
rect 4847 8585 4859 8588
rect 4801 8579 4859 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5353 8619 5411 8625
rect 5353 8585 5365 8619
rect 5399 8616 5411 8619
rect 5442 8616 5448 8628
rect 5399 8588 5448 8616
rect 5399 8585 5411 8588
rect 5353 8579 5411 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 6730 8616 6736 8628
rect 6687 8588 6736 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 7650 8616 7656 8628
rect 7423 8588 7656 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 8110 8616 8116 8628
rect 7791 8588 8116 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8478 8616 8484 8628
rect 8343 8588 8484 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8665 8619 8723 8625
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 8754 8616 8760 8628
rect 8711 8588 8760 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 9088 8588 9229 8616
rect 9088 8576 9094 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9217 8579 9275 8585
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9364 8588 9597 8616
rect 9364 8576 9370 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11480 8588 12081 8616
rect 11480 8576 11486 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 12069 8579 12127 8585
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 12345 8619 12403 8625
rect 12345 8616 12357 8619
rect 12216 8588 12357 8616
rect 12216 8576 12222 8588
rect 12345 8585 12357 8588
rect 12391 8585 12403 8619
rect 12345 8579 12403 8585
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 12676 8588 13093 8616
rect 12676 8576 12682 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 13906 8576 13912 8628
rect 13964 8576 13970 8628
rect 14182 8576 14188 8628
rect 14240 8616 14246 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 14240 8588 14381 8616
rect 14240 8576 14246 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 14369 8579 14427 8585
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14516 8588 14964 8616
rect 14516 8576 14522 8588
rect 716 8520 3188 8548
rect 3973 8551 4031 8557
rect 716 8508 722 8520
rect 3973 8517 3985 8551
rect 4019 8517 4031 8551
rect 3973 8511 4031 8517
rect 5077 8551 5135 8557
rect 5077 8517 5089 8551
rect 5123 8548 5135 8551
rect 7834 8548 7840 8560
rect 5123 8520 7840 8548
rect 5123 8517 5135 8520
rect 5077 8511 5135 8517
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 1964 8412 1992 8443
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2774 8480 2780 8492
rect 2746 8440 2780 8480
rect 2832 8440 2838 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 2746 8412 2774 8440
rect 1964 8384 2774 8412
rect 3068 8344 3096 8443
rect 3988 8412 4016 8511
rect 7834 8508 7840 8520
rect 7892 8508 7898 8560
rect 8018 8508 8024 8560
rect 8076 8508 8082 8560
rect 9950 8548 9956 8560
rect 8496 8520 9956 8548
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 5534 8480 5540 8492
rect 4663 8452 5540 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5626 8440 5632 8492
rect 5684 8440 5690 8492
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6638 8480 6644 8492
rect 6595 8452 6644 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8480 7251 8483
rect 7466 8480 7472 8492
rect 7239 8452 7472 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 8386 8480 8392 8492
rect 8128 8452 8392 8480
rect 8128 8412 8156 8452
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8496 8489 8524 8520
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 12636 8520 13860 8548
rect 12529 8492 12587 8493
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9214 8480 9220 8492
rect 9079 8452 9220 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 9398 8440 9404 8492
rect 9456 8440 9462 8492
rect 10042 8440 10048 8492
rect 10100 8440 10106 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10594 8480 10600 8492
rect 10275 8452 10600 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 11146 8480 11152 8492
rect 10735 8452 11152 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 11514 8480 11520 8492
rect 11379 8452 11520 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 9766 8412 9772 8424
rect 3988 8384 8156 8412
rect 8220 8384 9772 8412
rect 7466 8344 7472 8356
rect 3068 8316 7472 8344
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 8220 8344 8248 8384
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 9916 8384 10916 8412
rect 9916 8372 9922 8384
rect 7616 8316 8248 8344
rect 7616 8304 7622 8316
rect 9582 8304 9588 8356
rect 9640 8344 9646 8356
rect 10888 8353 10916 8384
rect 10980 8384 11652 8412
rect 10413 8347 10471 8353
rect 10413 8344 10425 8347
rect 9640 8316 10425 8344
rect 9640 8304 9646 8316
rect 10413 8313 10425 8316
rect 10459 8313 10471 8347
rect 10413 8307 10471 8313
rect 10873 8347 10931 8353
rect 10873 8313 10885 8347
rect 10919 8313 10931 8347
rect 10873 8307 10931 8313
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 8386 8276 8392 8288
rect 5960 8248 8392 8276
rect 5960 8236 5966 8248
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 9861 8279 9919 8285
rect 9861 8276 9873 8279
rect 8536 8248 9873 8276
rect 8536 8236 8542 8248
rect 9861 8245 9873 8248
rect 9907 8245 9919 8279
rect 9861 8239 9919 8245
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10980 8276 11008 8384
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11112 8316 11529 8344
rect 11112 8304 11118 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 10008 8248 11008 8276
rect 11149 8279 11207 8285
rect 10008 8236 10014 8248
rect 11149 8245 11161 8279
rect 11195 8276 11207 8279
rect 11330 8276 11336 8288
rect 11195 8248 11336 8276
rect 11195 8245 11207 8248
rect 11149 8239 11207 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11624 8276 11652 8384
rect 11716 8344 11744 8443
rect 11974 8440 11980 8492
rect 12032 8440 12038 8492
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12268 8412 12296 8443
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12636 8489 12664 8520
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12768 8452 12909 8480
rect 12768 8440 12774 8452
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13630 8440 13636 8492
rect 13688 8440 13694 8492
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 12434 8412 12440 8424
rect 12268 8384 12440 8412
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 12802 8372 12808 8424
rect 12860 8412 12866 8424
rect 12860 8384 13492 8412
rect 12860 8372 12866 8384
rect 13464 8353 13492 8384
rect 13173 8347 13231 8353
rect 13173 8344 13185 8347
rect 11716 8316 12388 8344
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 11624 8248 11805 8276
rect 11793 8245 11805 8248
rect 11839 8245 11851 8279
rect 12360 8276 12388 8316
rect 12544 8316 13185 8344
rect 12544 8276 12572 8316
rect 13173 8313 13185 8316
rect 13219 8313 13231 8347
rect 13173 8307 13231 8313
rect 13449 8347 13507 8353
rect 13449 8313 13461 8347
rect 13495 8313 13507 8347
rect 13449 8307 13507 8313
rect 12360 8248 12572 8276
rect 12805 8279 12863 8285
rect 11793 8239 11851 8245
rect 12805 8245 12817 8279
rect 12851 8276 12863 8279
rect 13556 8276 13584 8440
rect 13740 8344 13768 8443
rect 13832 8412 13860 8520
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 14056 8520 14688 8548
rect 14056 8508 14062 8520
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14458 8440 14464 8492
rect 14516 8440 14522 8492
rect 14660 8489 14688 8520
rect 14936 8489 14964 8588
rect 15194 8576 15200 8628
rect 15252 8576 15258 8628
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 15749 8619 15807 8625
rect 15749 8616 15761 8619
rect 15528 8588 15761 8616
rect 15528 8576 15534 8588
rect 15749 8585 15761 8588
rect 15795 8585 15807 8619
rect 15749 8579 15807 8585
rect 15838 8576 15844 8628
rect 15896 8576 15902 8628
rect 16117 8619 16175 8625
rect 16117 8585 16129 8619
rect 16163 8585 16175 8619
rect 16117 8579 16175 8585
rect 16132 8548 16160 8579
rect 16298 8576 16304 8628
rect 16356 8576 16362 8628
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 16448 8588 16528 8616
rect 16448 8576 16454 8588
rect 15580 8520 16160 8548
rect 16316 8548 16344 8576
rect 16500 8548 16528 8588
rect 16666 8576 16672 8628
rect 16724 8576 16730 8628
rect 16942 8576 16948 8628
rect 17000 8576 17006 8628
rect 17218 8576 17224 8628
rect 17276 8576 17282 8628
rect 17494 8576 17500 8628
rect 17552 8576 17558 8628
rect 17586 8576 17592 8628
rect 17644 8616 17650 8628
rect 17644 8588 18460 8616
rect 17644 8576 17650 8588
rect 16316 8520 16436 8548
rect 16500 8520 17908 8548
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 15194 8480 15200 8492
rect 15059 8452 15200 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 15580 8489 15608 8520
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8449 15623 8483
rect 15565 8443 15623 8449
rect 14476 8412 14504 8440
rect 13832 8384 14504 8412
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 15488 8412 15516 8443
rect 15654 8440 15660 8492
rect 15712 8480 15718 8492
rect 16025 8483 16083 8489
rect 16025 8480 16037 8483
rect 15712 8452 16037 8480
rect 15712 8440 15718 8452
rect 16025 8449 16037 8452
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8449 16359 8483
rect 16301 8443 16359 8449
rect 14608 8384 15516 8412
rect 14608 8372 14614 8384
rect 14366 8344 14372 8356
rect 13740 8316 14372 8344
rect 14366 8304 14372 8316
rect 14424 8304 14430 8356
rect 14458 8304 14464 8356
rect 14516 8304 14522 8356
rect 15289 8347 15347 8353
rect 15289 8344 15301 8347
rect 14568 8316 15301 8344
rect 14568 8288 14596 8316
rect 15289 8313 15301 8316
rect 15335 8313 15347 8347
rect 15289 8307 15347 8313
rect 15378 8304 15384 8356
rect 15436 8344 15442 8356
rect 16316 8344 16344 8443
rect 15436 8316 16344 8344
rect 16408 8344 16436 8520
rect 16850 8440 16856 8492
rect 16908 8440 16914 8492
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 17144 8412 17172 8443
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 16724 8384 17172 8412
rect 16724 8372 16730 8384
rect 17218 8372 17224 8424
rect 17276 8412 17282 8424
rect 17696 8412 17724 8443
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 17276 8384 17724 8412
rect 17880 8412 17908 8520
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18432 8480 18460 8588
rect 18598 8576 18604 8628
rect 18656 8616 18662 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 18656 8588 19073 8616
rect 18656 8576 18662 8588
rect 19061 8585 19073 8588
rect 19107 8585 19119 8619
rect 19061 8579 19119 8585
rect 19978 8576 19984 8628
rect 20036 8576 20042 8628
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20349 8619 20407 8625
rect 20349 8616 20361 8619
rect 20128 8588 20361 8616
rect 20128 8576 20134 8588
rect 20349 8585 20361 8588
rect 20395 8585 20407 8619
rect 20349 8579 20407 8585
rect 20530 8576 20536 8628
rect 20588 8616 20594 8628
rect 20717 8619 20775 8625
rect 20717 8616 20729 8619
rect 20588 8588 20729 8616
rect 20588 8576 20594 8588
rect 20717 8585 20729 8588
rect 20763 8585 20775 8619
rect 20717 8579 20775 8585
rect 20898 8576 20904 8628
rect 20956 8616 20962 8628
rect 21269 8619 21327 8625
rect 21269 8616 21281 8619
rect 20956 8588 21281 8616
rect 20956 8576 20962 8588
rect 21269 8585 21281 8588
rect 21315 8585 21327 8619
rect 21269 8579 21327 8585
rect 21542 8576 21548 8628
rect 21600 8616 21606 8628
rect 22373 8619 22431 8625
rect 22373 8616 22385 8619
rect 21600 8588 22385 8616
rect 21600 8576 21606 8588
rect 22373 8585 22385 8588
rect 22419 8585 22431 8619
rect 22373 8579 22431 8585
rect 22922 8576 22928 8628
rect 22980 8576 22986 8628
rect 23106 8576 23112 8628
rect 23164 8616 23170 8628
rect 23477 8619 23535 8625
rect 23477 8616 23489 8619
rect 23164 8588 23489 8616
rect 23164 8576 23170 8588
rect 23477 8585 23489 8588
rect 23523 8585 23535 8619
rect 23477 8579 23535 8585
rect 18966 8548 18972 8560
rect 18800 8520 18972 8548
rect 18800 8489 18828 8520
rect 18966 8508 18972 8520
rect 19024 8508 19030 8560
rect 19150 8508 19156 8560
rect 19208 8548 19214 8560
rect 19208 8520 19840 8548
rect 19208 8508 19214 8520
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18095 8452 18368 8480
rect 18432 8452 18521 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 17880 8384 18184 8412
rect 17276 8372 17282 8384
rect 17957 8347 18015 8353
rect 17957 8344 17969 8347
rect 16408 8316 17969 8344
rect 15436 8304 15442 8316
rect 17957 8313 17969 8316
rect 18003 8313 18015 8347
rect 17957 8307 18015 8313
rect 12851 8248 13584 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 14550 8236 14556 8288
rect 14608 8236 14614 8288
rect 14734 8236 14740 8288
rect 14792 8236 14798 8288
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 17862 8276 17868 8288
rect 15068 8248 17868 8276
rect 15068 8236 15074 8248
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 18156 8276 18184 8384
rect 18230 8304 18236 8356
rect 18288 8304 18294 8356
rect 18340 8353 18368 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 18598 8372 18604 8424
rect 18656 8412 18662 8424
rect 19444 8412 19472 8443
rect 19702 8440 19708 8492
rect 19760 8440 19766 8492
rect 19812 8489 19840 8520
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 20162 8440 20168 8492
rect 20220 8440 20226 8492
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8449 20683 8483
rect 20625 8443 20683 8449
rect 18656 8384 19472 8412
rect 18656 8372 18662 8384
rect 18325 8347 18383 8353
rect 18325 8313 18337 8347
rect 18371 8313 18383 8347
rect 20640 8344 20668 8443
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 21177 8483 21235 8489
rect 21177 8480 21189 8483
rect 20864 8452 21189 8480
rect 20864 8440 20870 8452
rect 21177 8449 21189 8452
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 21266 8440 21272 8492
rect 21324 8480 21330 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21324 8452 21833 8480
rect 21324 8440 21330 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22278 8440 22284 8492
rect 22336 8440 22342 8492
rect 22462 8440 22468 8492
rect 22520 8480 22526 8492
rect 22833 8483 22891 8489
rect 22833 8480 22845 8483
rect 22520 8452 22845 8480
rect 22520 8440 22526 8452
rect 22833 8449 22845 8452
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 22922 8440 22928 8492
rect 22980 8480 22986 8492
rect 23385 8483 23443 8489
rect 23385 8480 23397 8483
rect 22980 8452 23397 8480
rect 22980 8440 22986 8452
rect 23385 8449 23397 8452
rect 23431 8449 23443 8483
rect 23385 8443 23443 8449
rect 20990 8372 20996 8424
rect 21048 8372 21054 8424
rect 18325 8307 18383 8313
rect 18432 8316 20668 8344
rect 21008 8344 21036 8372
rect 22005 8347 22063 8353
rect 22005 8344 22017 8347
rect 21008 8316 22017 8344
rect 18432 8276 18460 8316
rect 22005 8313 22017 8316
rect 22051 8313 22063 8347
rect 22005 8307 22063 8313
rect 18156 8248 18460 8276
rect 18598 8236 18604 8288
rect 18656 8236 18662 8288
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 19245 8279 19303 8285
rect 19245 8276 19257 8279
rect 19208 8248 19257 8276
rect 19208 8236 19214 8248
rect 19245 8245 19257 8248
rect 19291 8245 19303 8279
rect 19245 8239 19303 8245
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 19521 8279 19579 8285
rect 19521 8276 19533 8279
rect 19392 8248 19533 8276
rect 19392 8236 19398 8248
rect 19521 8245 19533 8248
rect 19567 8245 19579 8279
rect 19521 8239 19579 8245
rect 1104 8186 24840 8208
rect 1104 8134 3917 8186
rect 3969 8134 3981 8186
rect 4033 8134 4045 8186
rect 4097 8134 4109 8186
rect 4161 8134 4173 8186
rect 4225 8134 9851 8186
rect 9903 8134 9915 8186
rect 9967 8134 9979 8186
rect 10031 8134 10043 8186
rect 10095 8134 10107 8186
rect 10159 8134 15785 8186
rect 15837 8134 15849 8186
rect 15901 8134 15913 8186
rect 15965 8134 15977 8186
rect 16029 8134 16041 8186
rect 16093 8134 21719 8186
rect 21771 8134 21783 8186
rect 21835 8134 21847 8186
rect 21899 8134 21911 8186
rect 21963 8134 21975 8186
rect 22027 8134 24840 8186
rect 1104 8112 24840 8134
rect 1670 8032 1676 8084
rect 1728 8032 1734 8084
rect 2406 8032 2412 8084
rect 2464 8032 2470 8084
rect 2774 8032 2780 8084
rect 2832 8032 2838 8084
rect 3326 8032 3332 8084
rect 3384 8032 3390 8084
rect 4154 8032 4160 8084
rect 4212 8032 4218 8084
rect 4982 8032 4988 8084
rect 5040 8032 5046 8084
rect 5902 8072 5908 8084
rect 5276 8044 5908 8072
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1762 7868 1768 7880
rect 1627 7840 1768 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7868 2191 7871
rect 2314 7868 2320 7880
rect 2179 7840 2320 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 3142 7868 3148 7880
rect 2731 7840 3148 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 5276 7868 5304 8044
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 6086 8032 6092 8084
rect 6144 8032 6150 8084
rect 6270 8032 6276 8084
rect 6328 8032 6334 8084
rect 6638 8032 6644 8084
rect 6696 8032 6702 8084
rect 7190 8032 7196 8084
rect 7248 8032 7254 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7432 8044 7757 8072
rect 7432 8032 7438 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8294 8032 8300 8084
rect 8352 8032 8358 8084
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 11057 8075 11115 8081
rect 11057 8072 11069 8075
rect 8444 8044 11069 8072
rect 8444 8032 8450 8044
rect 11057 8041 11069 8044
rect 11103 8041 11115 8075
rect 11057 8035 11115 8041
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 11204 8044 11621 8072
rect 11204 8032 11210 8044
rect 11609 8041 11621 8044
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 12176 8044 12572 8072
rect 5721 8007 5779 8013
rect 5721 7973 5733 8007
rect 5767 8004 5779 8007
rect 6288 8004 6316 8032
rect 9401 8007 9459 8013
rect 9401 8004 9413 8007
rect 5767 7976 6316 8004
rect 6748 7976 9413 8004
rect 5767 7973 5779 7976
rect 5721 7967 5779 7973
rect 5350 7896 5356 7948
rect 5408 7936 5414 7948
rect 6748 7936 6776 7976
rect 9401 7973 9413 7976
rect 9447 7973 9459 8007
rect 9401 7967 9459 7973
rect 9674 7964 9680 8016
rect 9732 7964 9738 8016
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 7973 9919 8007
rect 10870 8004 10876 8016
rect 9861 7967 9919 7973
rect 9968 7976 10876 8004
rect 7926 7936 7932 7948
rect 5408 7908 6776 7936
rect 7576 7908 7932 7936
rect 5408 7896 5414 7908
rect 4111 7840 5304 7868
rect 5537 7871 5595 7877
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 5810 7868 5816 7880
rect 5583 7840 5816 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 3252 7744 3280 7831
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 7576 7877 7604 7908
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 8628 7908 9260 7936
rect 8628 7896 8634 7908
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8938 7868 8944 7880
rect 8251 7840 8944 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7769 4951 7803
rect 4893 7763 4951 7769
rect 3234 7692 3240 7744
rect 3292 7692 3298 7744
rect 4908 7732 4936 7763
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 5997 7803 6055 7809
rect 5997 7800 6009 7803
rect 5500 7772 6009 7800
rect 5500 7760 5506 7772
rect 5997 7769 6009 7772
rect 6043 7769 6055 7803
rect 5997 7763 6055 7769
rect 6546 7760 6552 7812
rect 6604 7760 6610 7812
rect 7101 7803 7159 7809
rect 7101 7769 7113 7803
rect 7147 7800 7159 7803
rect 8110 7800 8116 7812
rect 7147 7772 8116 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 4908 7704 9137 7732
rect 9125 7701 9137 7704
rect 9171 7701 9183 7735
rect 9232 7732 9260 7908
rect 9692 7893 9720 7964
rect 9677 7887 9735 7893
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9324 7800 9352 7831
rect 9582 7828 9588 7880
rect 9640 7828 9646 7880
rect 9677 7853 9689 7887
rect 9723 7853 9735 7887
rect 9677 7847 9735 7853
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 9876 7868 9904 7967
rect 9824 7840 9904 7868
rect 9824 7828 9830 7840
rect 9968 7800 9996 7976
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 11333 8007 11391 8013
rect 11333 7973 11345 8007
rect 11379 7973 11391 8007
rect 11333 7967 11391 7973
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 11348 7936 11376 7967
rect 11514 7964 11520 8016
rect 11572 8004 11578 8016
rect 12176 8004 12204 8044
rect 12437 8007 12495 8013
rect 12437 8004 12449 8007
rect 11572 7976 12204 8004
rect 12268 7976 12449 8004
rect 11572 7964 11578 7976
rect 12158 7936 12164 7948
rect 10652 7908 11376 7936
rect 11440 7908 12164 7936
rect 10652 7896 10658 7908
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 9324 7772 9996 7800
rect 10152 7800 10180 7831
rect 10410 7828 10416 7880
rect 10468 7828 10474 7880
rect 10686 7828 10692 7880
rect 10744 7828 10750 7880
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7868 11299 7871
rect 11440 7868 11468 7908
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 11287 7840 11468 7868
rect 11287 7837 11299 7840
rect 11241 7831 11299 7837
rect 11514 7828 11520 7880
rect 11572 7828 11578 7880
rect 11790 7828 11796 7880
rect 11848 7828 11854 7880
rect 12066 7828 12072 7880
rect 12124 7828 12130 7880
rect 12268 7800 12296 7976
rect 12437 7973 12449 7976
rect 12483 7973 12495 8007
rect 12544 8004 12572 8044
rect 12986 8032 12992 8084
rect 13044 8032 13050 8084
rect 14090 8032 14096 8084
rect 14148 8032 14154 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14921 8075 14979 8081
rect 14921 8072 14933 8075
rect 14240 8044 14933 8072
rect 14240 8032 14246 8044
rect 14921 8041 14933 8044
rect 14967 8041 14979 8075
rect 14921 8035 14979 8041
rect 15194 8032 15200 8084
rect 15252 8032 15258 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 15841 8075 15899 8081
rect 15841 8072 15853 8075
rect 15712 8044 15853 8072
rect 15712 8032 15718 8044
rect 15841 8041 15853 8044
rect 15887 8041 15899 8075
rect 15841 8035 15899 8041
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16850 8072 16856 8084
rect 16439 8044 16856 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17402 8072 17408 8084
rect 16991 8044 17408 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8072 17555 8075
rect 17770 8072 17776 8084
rect 17543 8044 17776 8072
rect 17543 8041 17555 8044
rect 17497 8035 17555 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 17862 8032 17868 8084
rect 17920 8072 17926 8084
rect 17957 8075 18015 8081
rect 17957 8072 17969 8075
rect 17920 8044 17969 8072
rect 17920 8032 17926 8044
rect 17957 8041 17969 8044
rect 18003 8041 18015 8075
rect 18598 8072 18604 8084
rect 17957 8035 18015 8041
rect 18064 8044 18604 8072
rect 13265 8007 13323 8013
rect 13265 8004 13277 8007
rect 12544 7976 13277 8004
rect 12437 7967 12495 7973
rect 13265 7973 13277 7976
rect 13311 7973 13323 8007
rect 14108 8004 14136 8032
rect 15565 8007 15623 8013
rect 15565 8004 15577 8007
rect 14108 7976 15577 8004
rect 13265 7967 13323 7973
rect 15565 7973 15577 7976
rect 15611 7973 15623 8007
rect 15565 7967 15623 7973
rect 16117 8007 16175 8013
rect 16117 7973 16129 8007
rect 16163 7973 16175 8007
rect 16117 7967 16175 7973
rect 16132 7936 16160 7967
rect 16482 7964 16488 8016
rect 16540 8004 16546 8016
rect 16540 7976 16896 8004
rect 16540 7964 16546 7976
rect 15764 7908 16160 7936
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 12400 7840 12633 7868
rect 12400 7828 12406 7840
rect 12621 7837 12633 7840
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14884 7840 15117 7868
rect 14884 7828 14890 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15378 7828 15384 7880
rect 15436 7828 15442 7880
rect 15764 7877 15792 7908
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16264 7908 16620 7936
rect 16264 7896 16270 7908
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 10152 7772 12296 7800
rect 15654 7760 15660 7812
rect 15712 7800 15718 7812
rect 16040 7800 16068 7831
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 16592 7877 16620 7908
rect 16868 7877 16896 7976
rect 17218 7964 17224 8016
rect 17276 7964 17282 8016
rect 17310 7964 17316 8016
rect 17368 8004 17374 8016
rect 17368 7976 17724 8004
rect 17368 7964 17374 7976
rect 17034 7896 17040 7948
rect 17092 7936 17098 7948
rect 17092 7908 17448 7936
rect 17092 7896 17098 7908
rect 17420 7877 17448 7908
rect 17696 7877 17724 7976
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 16172 7840 16313 7868
rect 16172 7828 16178 7840
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 16853 7871 16911 7877
rect 16853 7837 16865 7871
rect 16899 7837 16911 7871
rect 16853 7831 16911 7837
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7868 17831 7871
rect 18064 7868 18092 8044
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 18874 8072 18880 8084
rect 18708 8044 18880 8072
rect 18233 8007 18291 8013
rect 18233 7973 18245 8007
rect 18279 8004 18291 8007
rect 18708 8004 18736 8044
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 19334 8032 19340 8084
rect 19392 8032 19398 8084
rect 21085 8075 21143 8081
rect 21085 8041 21097 8075
rect 21131 8072 21143 8075
rect 21174 8072 21180 8084
rect 21131 8044 21180 8072
rect 21131 8041 21143 8044
rect 21085 8035 21143 8041
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 22554 8032 22560 8084
rect 22612 8032 22618 8084
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 23109 8075 23167 8081
rect 23109 8072 23121 8075
rect 22888 8044 23121 8072
rect 22888 8032 22894 8044
rect 23109 8041 23121 8044
rect 23155 8041 23167 8075
rect 23109 8035 23167 8041
rect 23382 8032 23388 8084
rect 23440 8032 23446 8084
rect 23658 8032 23664 8084
rect 23716 8072 23722 8084
rect 23937 8075 23995 8081
rect 23937 8072 23949 8075
rect 23716 8044 23949 8072
rect 23716 8032 23722 8044
rect 23937 8041 23949 8044
rect 23983 8041 23995 8075
rect 23937 8035 23995 8041
rect 18279 7976 18736 8004
rect 18279 7973 18291 7976
rect 18233 7967 18291 7973
rect 18782 7964 18788 8016
rect 18840 8004 18846 8016
rect 18969 8007 19027 8013
rect 18969 8004 18981 8007
rect 18840 7976 18981 8004
rect 18840 7964 18846 7976
rect 18969 7973 18981 7976
rect 19015 7973 19027 8007
rect 18969 7967 19027 7973
rect 19352 7936 19380 8032
rect 22189 8007 22247 8013
rect 22189 7973 22201 8007
rect 22235 8004 22247 8007
rect 23400 8004 23428 8032
rect 22235 7976 23428 8004
rect 22235 7973 22247 7976
rect 22189 7967 22247 7973
rect 18800 7908 19380 7936
rect 17819 7840 18092 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 15712 7772 16068 7800
rect 15712 7760 15718 7772
rect 16758 7760 16764 7812
rect 16816 7800 16822 7812
rect 17144 7800 17172 7831
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18800 7877 18828 7908
rect 18417 7871 18475 7877
rect 18417 7868 18429 7871
rect 18196 7840 18429 7868
rect 18196 7828 18202 7840
rect 18417 7837 18429 7840
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7837 18843 7871
rect 18785 7831 18843 7837
rect 16816 7772 17172 7800
rect 18524 7800 18552 7831
rect 19150 7828 19156 7880
rect 19208 7828 19214 7880
rect 19334 7828 19340 7880
rect 19392 7828 19398 7880
rect 19610 7828 19616 7880
rect 19668 7828 19674 7880
rect 19886 7828 19892 7880
rect 19944 7828 19950 7880
rect 20898 7828 20904 7880
rect 20956 7828 20962 7880
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7868 21787 7871
rect 25590 7868 25596 7880
rect 21775 7840 25596 7868
rect 21775 7837 21787 7840
rect 21729 7831 21787 7837
rect 25590 7828 25596 7840
rect 25648 7828 25654 7880
rect 19168 7800 19196 7828
rect 18524 7772 19196 7800
rect 21361 7803 21419 7809
rect 16816 7760 16822 7772
rect 21361 7769 21373 7803
rect 21407 7800 21419 7803
rect 21407 7772 21772 7800
rect 21407 7769 21419 7772
rect 21361 7763 21419 7769
rect 9953 7735 10011 7741
rect 9953 7732 9965 7735
rect 9232 7704 9965 7732
rect 9125 7695 9183 7701
rect 9953 7701 9965 7704
rect 9999 7701 10011 7735
rect 9953 7695 10011 7701
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10229 7735 10287 7741
rect 10229 7732 10241 7735
rect 10100 7704 10241 7732
rect 10100 7692 10106 7704
rect 10229 7701 10241 7704
rect 10275 7701 10287 7735
rect 10229 7695 10287 7701
rect 10502 7692 10508 7744
rect 10560 7692 10566 7744
rect 10778 7692 10784 7744
rect 10836 7692 10842 7744
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11885 7735 11943 7741
rect 11885 7732 11897 7735
rect 10928 7704 11897 7732
rect 10928 7692 10934 7704
rect 11885 7701 11897 7704
rect 11931 7701 11943 7735
rect 11885 7695 11943 7701
rect 16666 7692 16672 7744
rect 16724 7692 16730 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 18693 7735 18751 7741
rect 18693 7732 18705 7735
rect 18104 7704 18705 7732
rect 18104 7692 18110 7704
rect 18693 7701 18705 7704
rect 18739 7701 18751 7735
rect 18693 7695 18751 7701
rect 19518 7692 19524 7744
rect 19576 7692 19582 7744
rect 19794 7692 19800 7744
rect 19852 7692 19858 7744
rect 20070 7692 20076 7744
rect 20128 7692 20134 7744
rect 21744 7732 21772 7772
rect 21910 7760 21916 7812
rect 21968 7760 21974 7812
rect 22462 7760 22468 7812
rect 22520 7760 22526 7812
rect 22646 7760 22652 7812
rect 22704 7800 22710 7812
rect 23017 7803 23075 7809
rect 23017 7800 23029 7803
rect 22704 7772 23029 7800
rect 22704 7760 22710 7772
rect 23017 7769 23029 7772
rect 23063 7769 23075 7803
rect 23017 7763 23075 7769
rect 23842 7760 23848 7812
rect 23900 7760 23906 7812
rect 23750 7732 23756 7744
rect 21744 7704 23756 7732
rect 23750 7692 23756 7704
rect 23808 7692 23814 7744
rect 1104 7642 25000 7664
rect 1104 7590 6884 7642
rect 6936 7590 6948 7642
rect 7000 7590 7012 7642
rect 7064 7590 7076 7642
rect 7128 7590 7140 7642
rect 7192 7590 12818 7642
rect 12870 7590 12882 7642
rect 12934 7590 12946 7642
rect 12998 7590 13010 7642
rect 13062 7590 13074 7642
rect 13126 7590 18752 7642
rect 18804 7590 18816 7642
rect 18868 7590 18880 7642
rect 18932 7590 18944 7642
rect 18996 7590 19008 7642
rect 19060 7590 24686 7642
rect 24738 7590 24750 7642
rect 24802 7590 24814 7642
rect 24866 7590 24878 7642
rect 24930 7590 24942 7642
rect 24994 7590 25000 7642
rect 1104 7568 25000 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 2041 7531 2099 7537
rect 2041 7528 2053 7531
rect 1360 7500 2053 7528
rect 1360 7488 1366 7500
rect 2041 7497 2053 7500
rect 2087 7497 2099 7531
rect 2041 7491 2099 7497
rect 2222 7488 2228 7540
rect 2280 7528 2286 7540
rect 2777 7531 2835 7537
rect 2777 7528 2789 7531
rect 2280 7500 2789 7528
rect 2280 7488 2286 7500
rect 2777 7497 2789 7500
rect 2823 7497 2835 7531
rect 2777 7491 2835 7497
rect 3513 7531 3571 7537
rect 3513 7497 3525 7531
rect 3559 7528 3571 7531
rect 3786 7528 3792 7540
rect 3559 7500 3792 7528
rect 3559 7497 3571 7500
rect 3513 7491 3571 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 4614 7488 4620 7540
rect 4672 7488 4678 7540
rect 5350 7488 5356 7540
rect 5408 7488 5414 7540
rect 5442 7488 5448 7540
rect 5500 7488 5506 7540
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 5684 7500 5733 7528
rect 5684 7488 5690 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 5997 7531 6055 7537
rect 5997 7528 6009 7531
rect 5868 7500 6009 7528
rect 5868 7488 5874 7500
rect 5997 7497 6009 7500
rect 6043 7497 6055 7531
rect 5997 7491 6055 7497
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6604 7500 6653 7528
rect 6604 7488 6610 7500
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 6641 7491 6699 7497
rect 7466 7488 7472 7540
rect 7524 7488 7530 7540
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7892 7500 8033 7528
rect 7892 7488 7898 7500
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 8021 7491 8079 7497
rect 8573 7531 8631 7537
rect 8573 7497 8585 7531
rect 8619 7528 8631 7531
rect 8662 7528 8668 7540
rect 8619 7500 8668 7528
rect 8619 7497 8631 7500
rect 8573 7491 8631 7497
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 10229 7531 10287 7537
rect 10229 7528 10241 7531
rect 9732 7500 10241 7528
rect 9732 7488 9738 7500
rect 10229 7497 10241 7500
rect 10275 7497 10287 7531
rect 10229 7491 10287 7497
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 11146 7528 11152 7540
rect 10376 7500 11152 7528
rect 10376 7488 10382 7500
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 21910 7528 21916 7540
rect 17828 7500 21916 7528
rect 17828 7488 17834 7500
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 22281 7531 22339 7537
rect 22281 7497 22293 7531
rect 22327 7528 22339 7531
rect 22554 7528 22560 7540
rect 22327 7500 22560 7528
rect 22327 7497 22339 7500
rect 22281 7491 22339 7497
rect 22554 7488 22560 7500
rect 22612 7488 22618 7540
rect 23937 7531 23995 7537
rect 23937 7497 23949 7531
rect 23983 7528 23995 7531
rect 24210 7528 24216 7540
rect 23983 7500 24216 7528
rect 23983 7497 23995 7500
rect 23937 7491 23995 7497
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 25314 7488 25320 7540
rect 25372 7488 25378 7540
rect 1946 7420 1952 7472
rect 2004 7420 2010 7472
rect 2501 7463 2559 7469
rect 2501 7429 2513 7463
rect 2547 7460 2559 7463
rect 2682 7460 2688 7472
rect 2547 7432 2688 7460
rect 2547 7429 2559 7432
rect 2501 7423 2559 7429
rect 2682 7420 2688 7432
rect 2740 7420 2746 7472
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7392 3387 7395
rect 4433 7395 4491 7401
rect 3375 7364 4384 7392
rect 3375 7361 3387 7364
rect 3329 7355 3387 7361
rect 2976 7324 3004 7355
rect 2976 7296 3648 7324
rect 3145 7191 3203 7197
rect 3145 7157 3157 7191
rect 3191 7188 3203 7191
rect 3510 7188 3516 7200
rect 3191 7160 3516 7188
rect 3191 7157 3203 7160
rect 3145 7151 3203 7157
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 3620 7188 3648 7296
rect 4356 7256 4384 7364
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 5368 7392 5396 7488
rect 19794 7460 19800 7472
rect 5644 7432 19800 7460
rect 5644 7401 5672 7432
rect 19794 7420 19800 7432
rect 19852 7420 19858 7472
rect 22925 7463 22983 7469
rect 22925 7429 22937 7463
rect 22971 7460 22983 7463
rect 25332 7460 25360 7488
rect 22971 7432 25360 7460
rect 22971 7429 22983 7432
rect 22925 7423 22983 7429
rect 4479 7364 5396 7392
rect 5629 7395 5687 7401
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 5629 7361 5641 7395
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 6871 7364 7205 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7193 7361 7205 7364
rect 7239 7392 7251 7395
rect 7558 7392 7564 7404
rect 7239 7364 7564 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 6564 7324 6592 7355
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8662 7392 8668 7404
rect 8251 7364 8668 7392
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 7374 7324 7380 7336
rect 6564 7296 7380 7324
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7668 7256 7696 7355
rect 7944 7324 7972 7355
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 10318 7392 10324 7404
rect 8803 7364 10324 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 10778 7352 10784 7404
rect 10836 7352 10842 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 20772 7364 22017 7392
rect 20772 7352 20778 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 10796 7324 10824 7352
rect 7944 7296 10824 7324
rect 22572 7324 22600 7355
rect 23106 7352 23112 7404
rect 23164 7352 23170 7404
rect 23658 7352 23664 7404
rect 23716 7352 23722 7404
rect 23290 7324 23296 7336
rect 22572 7296 23296 7324
rect 23290 7284 23296 7296
rect 23348 7284 23354 7336
rect 23385 7327 23443 7333
rect 23385 7293 23397 7327
rect 23431 7324 23443 7327
rect 25038 7324 25044 7336
rect 23431 7296 25044 7324
rect 23431 7293 23443 7296
rect 23385 7287 23443 7293
rect 25038 7284 25044 7296
rect 25096 7284 25102 7336
rect 10502 7256 10508 7268
rect 4356 7228 7236 7256
rect 7668 7228 10508 7256
rect 6270 7188 6276 7200
rect 3620 7160 6276 7188
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6362 7148 6368 7200
rect 6420 7148 6426 7200
rect 7208 7188 7236 7228
rect 10502 7216 10508 7228
rect 10560 7216 10566 7268
rect 10594 7216 10600 7268
rect 10652 7216 10658 7268
rect 8478 7188 8484 7200
rect 7208 7160 8484 7188
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 10612 7188 10640 7216
rect 8720 7160 10640 7188
rect 8720 7148 8726 7160
rect 1104 7098 24840 7120
rect 1104 7046 3917 7098
rect 3969 7046 3981 7098
rect 4033 7046 4045 7098
rect 4097 7046 4109 7098
rect 4161 7046 4173 7098
rect 4225 7046 9851 7098
rect 9903 7046 9915 7098
rect 9967 7046 9979 7098
rect 10031 7046 10043 7098
rect 10095 7046 10107 7098
rect 10159 7046 15785 7098
rect 15837 7046 15849 7098
rect 15901 7046 15913 7098
rect 15965 7046 15977 7098
rect 16029 7046 16041 7098
rect 16093 7046 21719 7098
rect 21771 7046 21783 7098
rect 21835 7046 21847 7098
rect 21899 7046 21911 7098
rect 21963 7046 21975 7098
rect 22027 7046 24840 7098
rect 1104 7024 24840 7046
rect 3234 6944 3240 6996
rect 3292 6984 3298 6996
rect 11054 6984 11060 6996
rect 3292 6956 11060 6984
rect 3292 6944 3298 6956
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 11330 6944 11336 6996
rect 11388 6944 11394 6996
rect 18046 6984 18052 6996
rect 12406 6956 18052 6984
rect 6270 6876 6276 6928
rect 6328 6916 6334 6928
rect 11348 6916 11376 6944
rect 6328 6888 11376 6916
rect 6328 6876 6334 6888
rect 1026 6808 1032 6860
rect 1084 6848 1090 6860
rect 1949 6851 2007 6857
rect 1949 6848 1961 6851
rect 1084 6820 1961 6848
rect 1084 6808 1090 6820
rect 1949 6817 1961 6820
rect 1995 6817 2007 6851
rect 1949 6811 2007 6817
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 12406 6848 12434 6956
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 22094 6944 22100 6996
rect 22152 6984 22158 6996
rect 23109 6987 23167 6993
rect 23109 6984 23121 6987
rect 22152 6956 23121 6984
rect 22152 6944 22158 6956
rect 23109 6953 23121 6956
rect 23155 6953 23167 6987
rect 23109 6947 23167 6953
rect 8168 6820 12434 6848
rect 23937 6851 23995 6857
rect 8168 6808 8174 6820
rect 23937 6817 23949 6851
rect 23983 6848 23995 6851
rect 24578 6848 24584 6860
rect 23983 6820 24584 6848
rect 23983 6817 23995 6820
rect 23937 6811 23995 6817
rect 24578 6808 24584 6820
rect 24636 6808 24642 6860
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 9766 6780 9772 6792
rect 1719 6752 9772 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 22094 6740 22100 6792
rect 22152 6780 22158 6792
rect 23661 6783 23719 6789
rect 23661 6780 23673 6783
rect 22152 6752 23673 6780
rect 22152 6740 22158 6752
rect 23661 6749 23673 6752
rect 23707 6749 23719 6783
rect 23661 6743 23719 6749
rect 2225 6715 2283 6721
rect 2225 6681 2237 6715
rect 2271 6712 2283 6715
rect 7742 6712 7748 6724
rect 2271 6684 7748 6712
rect 2271 6681 2283 6684
rect 2225 6675 2283 6681
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 23014 6672 23020 6724
rect 23072 6672 23078 6724
rect 198 6604 204 6656
rect 256 6644 262 6656
rect 2317 6647 2375 6653
rect 2317 6644 2329 6647
rect 256 6616 2329 6644
rect 256 6604 262 6616
rect 2317 6613 2329 6616
rect 2363 6613 2375 6647
rect 2317 6607 2375 6613
rect 1104 6554 25000 6576
rect 1104 6502 6884 6554
rect 6936 6502 6948 6554
rect 7000 6502 7012 6554
rect 7064 6502 7076 6554
rect 7128 6502 7140 6554
rect 7192 6502 12818 6554
rect 12870 6502 12882 6554
rect 12934 6502 12946 6554
rect 12998 6502 13010 6554
rect 13062 6502 13074 6554
rect 13126 6502 18752 6554
rect 18804 6502 18816 6554
rect 18868 6502 18880 6554
rect 18932 6502 18944 6554
rect 18996 6502 19008 6554
rect 19060 6502 24686 6554
rect 24738 6502 24750 6554
rect 24802 6502 24814 6554
rect 24866 6502 24878 6554
rect 24930 6502 24942 6554
rect 24994 6502 25000 6554
rect 1104 6480 25000 6502
rect 750 6400 756 6452
rect 808 6440 814 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 808 6412 1593 6440
rect 808 6400 814 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 23753 6443 23811 6449
rect 23753 6409 23765 6443
rect 23799 6440 23811 6443
rect 23934 6440 23940 6452
rect 23799 6412 23940 6440
rect 23799 6409 23811 6412
rect 23753 6403 23811 6409
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 24305 6443 24363 6449
rect 24305 6409 24317 6443
rect 24351 6440 24363 6443
rect 24486 6440 24492 6452
rect 24351 6412 24492 6440
rect 24351 6409 24363 6412
rect 24305 6403 24363 6409
rect 24486 6400 24492 6412
rect 24544 6400 24550 6452
rect 1489 6375 1547 6381
rect 1489 6341 1501 6375
rect 1535 6372 1547 6375
rect 6362 6372 6368 6384
rect 1535 6344 6368 6372
rect 1535 6341 1547 6344
rect 1489 6335 1547 6341
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 23382 6332 23388 6384
rect 23440 6372 23446 6384
rect 24029 6375 24087 6381
rect 24029 6372 24041 6375
rect 23440 6344 24041 6372
rect 23440 6332 23446 6344
rect 24029 6341 24041 6344
rect 24075 6341 24087 6375
rect 24029 6335 24087 6341
rect 17494 6264 17500 6316
rect 17552 6264 17558 6316
rect 23474 6264 23480 6316
rect 23532 6264 23538 6316
rect 17313 6103 17371 6109
rect 17313 6069 17325 6103
rect 17359 6100 17371 6103
rect 23842 6100 23848 6112
rect 17359 6072 23848 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 23842 6060 23848 6072
rect 23900 6060 23906 6112
rect 1104 6010 24840 6032
rect 1104 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 9851 6010
rect 9903 5958 9915 6010
rect 9967 5958 9979 6010
rect 10031 5958 10043 6010
rect 10095 5958 10107 6010
rect 10159 5958 15785 6010
rect 15837 5958 15849 6010
rect 15901 5958 15913 6010
rect 15965 5958 15977 6010
rect 16029 5958 16041 6010
rect 16093 5958 21719 6010
rect 21771 5958 21783 6010
rect 21835 5958 21847 6010
rect 21899 5958 21911 6010
rect 21963 5958 21975 6010
rect 22027 5958 24840 6010
rect 1104 5936 24840 5958
rect 16761 5899 16819 5905
rect 16761 5865 16773 5899
rect 16807 5896 16819 5899
rect 17494 5896 17500 5908
rect 16807 5868 17500 5896
rect 16807 5865 16819 5868
rect 16761 5859 16819 5865
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 16942 5652 16948 5704
rect 17000 5652 17006 5704
rect 1104 5466 25000 5488
rect 1104 5414 6884 5466
rect 6936 5414 6948 5466
rect 7000 5414 7012 5466
rect 7064 5414 7076 5466
rect 7128 5414 7140 5466
rect 7192 5414 12818 5466
rect 12870 5414 12882 5466
rect 12934 5414 12946 5466
rect 12998 5414 13010 5466
rect 13062 5414 13074 5466
rect 13126 5414 18752 5466
rect 18804 5414 18816 5466
rect 18868 5414 18880 5466
rect 18932 5414 18944 5466
rect 18996 5414 19008 5466
rect 19060 5414 24686 5466
rect 24738 5414 24750 5466
rect 24802 5414 24814 5466
rect 24866 5414 24878 5466
rect 24930 5414 24942 5466
rect 24994 5414 25000 5466
rect 1104 5392 25000 5414
rect 1104 4922 24840 4944
rect 1104 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 9851 4922
rect 9903 4870 9915 4922
rect 9967 4870 9979 4922
rect 10031 4870 10043 4922
rect 10095 4870 10107 4922
rect 10159 4870 15785 4922
rect 15837 4870 15849 4922
rect 15901 4870 15913 4922
rect 15965 4870 15977 4922
rect 16029 4870 16041 4922
rect 16093 4870 21719 4922
rect 21771 4870 21783 4922
rect 21835 4870 21847 4922
rect 21899 4870 21911 4922
rect 21963 4870 21975 4922
rect 22027 4870 24840 4922
rect 1104 4848 24840 4870
rect 1104 4378 25000 4400
rect 1104 4326 6884 4378
rect 6936 4326 6948 4378
rect 7000 4326 7012 4378
rect 7064 4326 7076 4378
rect 7128 4326 7140 4378
rect 7192 4326 12818 4378
rect 12870 4326 12882 4378
rect 12934 4326 12946 4378
rect 12998 4326 13010 4378
rect 13062 4326 13074 4378
rect 13126 4326 18752 4378
rect 18804 4326 18816 4378
rect 18868 4326 18880 4378
rect 18932 4326 18944 4378
rect 18996 4326 19008 4378
rect 19060 4326 24686 4378
rect 24738 4326 24750 4378
rect 24802 4326 24814 4378
rect 24866 4326 24878 4378
rect 24930 4326 24942 4378
rect 24994 4326 25000 4378
rect 1104 4304 25000 4326
rect 1104 3834 24840 3856
rect 1104 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 9851 3834
rect 9903 3782 9915 3834
rect 9967 3782 9979 3834
rect 10031 3782 10043 3834
rect 10095 3782 10107 3834
rect 10159 3782 15785 3834
rect 15837 3782 15849 3834
rect 15901 3782 15913 3834
rect 15965 3782 15977 3834
rect 16029 3782 16041 3834
rect 16093 3782 21719 3834
rect 21771 3782 21783 3834
rect 21835 3782 21847 3834
rect 21899 3782 21911 3834
rect 21963 3782 21975 3834
rect 22027 3782 24840 3834
rect 1104 3760 24840 3782
rect 1104 3290 25000 3312
rect 1104 3238 6884 3290
rect 6936 3238 6948 3290
rect 7000 3238 7012 3290
rect 7064 3238 7076 3290
rect 7128 3238 7140 3290
rect 7192 3238 12818 3290
rect 12870 3238 12882 3290
rect 12934 3238 12946 3290
rect 12998 3238 13010 3290
rect 13062 3238 13074 3290
rect 13126 3238 18752 3290
rect 18804 3238 18816 3290
rect 18868 3238 18880 3290
rect 18932 3238 18944 3290
rect 18996 3238 19008 3290
rect 19060 3238 24686 3290
rect 24738 3238 24750 3290
rect 24802 3238 24814 3290
rect 24866 3238 24878 3290
rect 24930 3238 24942 3290
rect 24994 3238 25000 3290
rect 1104 3216 25000 3238
rect 1104 2746 24840 2768
rect 1104 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 9851 2746
rect 9903 2694 9915 2746
rect 9967 2694 9979 2746
rect 10031 2694 10043 2746
rect 10095 2694 10107 2746
rect 10159 2694 15785 2746
rect 15837 2694 15849 2746
rect 15901 2694 15913 2746
rect 15965 2694 15977 2746
rect 16029 2694 16041 2746
rect 16093 2694 21719 2746
rect 21771 2694 21783 2746
rect 21835 2694 21847 2746
rect 21899 2694 21911 2746
rect 21963 2694 21975 2746
rect 22027 2694 24840 2746
rect 1104 2672 24840 2694
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 22646 2632 22652 2644
rect 13872 2604 22652 2632
rect 13872 2592 13878 2604
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 22922 2592 22928 2644
rect 22980 2592 22986 2644
rect 15102 2524 15108 2576
rect 15160 2564 15166 2576
rect 22940 2564 22968 2592
rect 15160 2536 22968 2564
rect 15160 2524 15166 2536
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 21266 2428 21272 2440
rect 13780 2400 21272 2428
rect 13780 2388 13786 2400
rect 21266 2388 21272 2400
rect 21324 2388 21330 2440
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 23658 2428 23664 2440
rect 22428 2400 23664 2428
rect 22428 2388 22434 2400
rect 23658 2388 23664 2400
rect 23716 2388 23722 2440
rect 23290 2320 23296 2372
rect 23348 2360 23354 2372
rect 24118 2360 24124 2372
rect 23348 2332 24124 2360
rect 23348 2320 23354 2332
rect 24118 2320 24124 2332
rect 24176 2320 24182 2372
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 20898 2292 20904 2304
rect 10652 2264 20904 2292
rect 10652 2252 10658 2264
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 1104 2202 25000 2224
rect 1104 2150 6884 2202
rect 6936 2150 6948 2202
rect 7000 2150 7012 2202
rect 7064 2150 7076 2202
rect 7128 2150 7140 2202
rect 7192 2150 12818 2202
rect 12870 2150 12882 2202
rect 12934 2150 12946 2202
rect 12998 2150 13010 2202
rect 13062 2150 13074 2202
rect 13126 2150 18752 2202
rect 18804 2150 18816 2202
rect 18868 2150 18880 2202
rect 18932 2150 18944 2202
rect 18996 2150 19008 2202
rect 19060 2150 24686 2202
rect 24738 2150 24750 2202
rect 24802 2150 24814 2202
rect 24866 2150 24878 2202
rect 24930 2150 24942 2202
rect 24994 2150 25000 2202
rect 1104 2128 25000 2150
rect 9122 2048 9128 2100
rect 9180 2048 9186 2100
rect 10226 2048 10232 2100
rect 10284 2048 10290 2100
rect 10594 2048 10600 2100
rect 10652 2048 10658 2100
rect 11698 2048 11704 2100
rect 11756 2048 11762 2100
rect 12805 2091 12863 2097
rect 12805 2057 12817 2091
rect 12851 2057 12863 2091
rect 12805 2051 12863 2057
rect 13081 2091 13139 2097
rect 13081 2057 13093 2091
rect 13127 2088 13139 2091
rect 13722 2088 13728 2100
rect 13127 2060 13728 2088
rect 13127 2057 13139 2060
rect 13081 2051 13139 2057
rect 12820 2020 12848 2051
rect 13722 2048 13728 2060
rect 13780 2048 13786 2100
rect 13814 2048 13820 2100
rect 13872 2048 13878 2100
rect 15102 2048 15108 2100
rect 15160 2048 15166 2100
rect 16301 2091 16359 2097
rect 16301 2057 16313 2091
rect 16347 2088 16359 2091
rect 17770 2088 17776 2100
rect 16347 2060 17776 2088
rect 16347 2057 16359 2060
rect 16301 2051 16359 2057
rect 17770 2048 17776 2060
rect 17828 2048 17834 2100
rect 20349 2091 20407 2097
rect 20349 2057 20361 2091
rect 20395 2057 20407 2091
rect 20349 2051 20407 2057
rect 20364 2020 20392 2051
rect 22094 2048 22100 2100
rect 22152 2048 22158 2100
rect 22370 2048 22376 2100
rect 22428 2048 22434 2100
rect 23106 2048 23112 2100
rect 23164 2088 23170 2100
rect 23569 2091 23627 2097
rect 23569 2088 23581 2091
rect 23164 2060 23581 2088
rect 23164 2048 23170 2060
rect 23569 2057 23581 2060
rect 23615 2057 23627 2091
rect 23569 2051 23627 2057
rect 23750 2048 23756 2100
rect 23808 2088 23814 2100
rect 23845 2091 23903 2097
rect 23845 2088 23857 2091
rect 23808 2060 23857 2088
rect 23808 2048 23814 2060
rect 23845 2057 23857 2060
rect 23891 2057 23903 2091
rect 23845 2051 23903 2057
rect 24118 2048 24124 2100
rect 24176 2048 24182 2100
rect 12820 1992 16804 2020
rect 20364 1992 23520 2020
rect 7742 1912 7748 1964
rect 7800 1912 7806 1964
rect 8938 1912 8944 1964
rect 8996 1912 9002 1964
rect 9766 1912 9772 1964
rect 9824 1952 9830 1964
rect 10045 1955 10103 1961
rect 10045 1952 10057 1955
rect 9824 1924 10057 1952
rect 9824 1912 9830 1924
rect 10045 1921 10057 1924
rect 10091 1921 10103 1955
rect 10045 1915 10103 1921
rect 10410 1912 10416 1964
rect 10468 1912 10474 1964
rect 11514 1912 11520 1964
rect 11572 1912 11578 1964
rect 12618 1912 12624 1964
rect 12676 1912 12682 1964
rect 12894 1912 12900 1964
rect 12952 1912 12958 1964
rect 13630 1912 13636 1964
rect 13688 1912 13694 1964
rect 13906 1912 13912 1964
rect 13964 1912 13970 1964
rect 14918 1912 14924 1964
rect 14976 1912 14982 1964
rect 15378 1912 15384 1964
rect 15436 1912 15442 1964
rect 16114 1912 16120 1964
rect 16172 1912 16178 1964
rect 16298 1912 16304 1964
rect 16356 1912 16362 1964
rect 7926 1776 7932 1828
rect 7984 1776 7990 1828
rect 14093 1819 14151 1825
rect 14093 1785 14105 1819
rect 14139 1816 14151 1819
rect 16316 1816 16344 1912
rect 16776 1884 16804 1992
rect 18598 1912 18604 1964
rect 18656 1912 18662 1964
rect 20530 1912 20536 1964
rect 20588 1912 20594 1964
rect 20714 1912 20720 1964
rect 20772 1912 20778 1964
rect 22278 1912 22284 1964
rect 22336 1912 22342 1964
rect 22554 1912 22560 1964
rect 22612 1912 22618 1964
rect 23492 1961 23520 1992
rect 23477 1955 23535 1961
rect 23477 1921 23489 1955
rect 23523 1921 23535 1955
rect 23477 1915 23535 1921
rect 23566 1912 23572 1964
rect 23624 1952 23630 1964
rect 23753 1955 23811 1961
rect 23753 1952 23765 1955
rect 23624 1924 23765 1952
rect 23624 1912 23630 1924
rect 23753 1921 23765 1924
rect 23799 1921 23811 1955
rect 23753 1915 23811 1921
rect 24026 1912 24032 1964
rect 24084 1912 24090 1964
rect 24302 1912 24308 1964
rect 24360 1912 24366 1964
rect 20732 1884 20760 1912
rect 16776 1856 20760 1884
rect 22066 1856 23520 1884
rect 14139 1788 16344 1816
rect 18785 1819 18843 1825
rect 14139 1785 14151 1788
rect 14093 1779 14151 1785
rect 18785 1785 18797 1819
rect 18831 1816 18843 1819
rect 22066 1816 22094 1856
rect 23492 1828 23520 1856
rect 18831 1788 22094 1816
rect 18831 1785 18843 1788
rect 18785 1779 18843 1785
rect 23382 1776 23388 1828
rect 23440 1776 23446 1828
rect 23474 1776 23480 1828
rect 23532 1776 23538 1828
rect 15565 1751 15623 1757
rect 15565 1717 15577 1751
rect 15611 1748 15623 1751
rect 20806 1748 20812 1760
rect 15611 1720 20812 1748
rect 15611 1717 15623 1720
rect 15565 1711 15623 1717
rect 20806 1708 20812 1720
rect 20864 1708 20870 1760
rect 23293 1751 23351 1757
rect 23293 1717 23305 1751
rect 23339 1748 23351 1751
rect 23400 1748 23428 1776
rect 23339 1720 23428 1748
rect 23339 1717 23351 1720
rect 23293 1711 23351 1717
rect 1104 1658 24840 1680
rect 1104 1606 3917 1658
rect 3969 1606 3981 1658
rect 4033 1606 4045 1658
rect 4097 1606 4109 1658
rect 4161 1606 4173 1658
rect 4225 1606 9851 1658
rect 9903 1606 9915 1658
rect 9967 1606 9979 1658
rect 10031 1606 10043 1658
rect 10095 1606 10107 1658
rect 10159 1606 15785 1658
rect 15837 1606 15849 1658
rect 15901 1606 15913 1658
rect 15965 1606 15977 1658
rect 16029 1606 16041 1658
rect 16093 1606 21719 1658
rect 21771 1606 21783 1658
rect 21835 1606 21847 1658
rect 21899 1606 21911 1658
rect 21963 1606 21975 1658
rect 22027 1606 24840 1658
rect 1104 1584 24840 1606
rect 7193 1547 7251 1553
rect 7193 1513 7205 1547
rect 7239 1544 7251 1547
rect 7742 1544 7748 1556
rect 7239 1516 7748 1544
rect 7239 1513 7251 1516
rect 7193 1507 7251 1513
rect 7742 1504 7748 1516
rect 7800 1504 7806 1556
rect 8389 1547 8447 1553
rect 8389 1513 8401 1547
rect 8435 1544 8447 1547
rect 8938 1544 8944 1556
rect 8435 1516 8944 1544
rect 8435 1513 8447 1516
rect 8389 1507 8447 1513
rect 8938 1504 8944 1516
rect 8996 1504 9002 1556
rect 9585 1547 9643 1553
rect 9585 1513 9597 1547
rect 9631 1544 9643 1547
rect 9766 1544 9772 1556
rect 9631 1516 9772 1544
rect 9631 1513 9643 1516
rect 9585 1507 9643 1513
rect 9766 1504 9772 1516
rect 9824 1504 9830 1556
rect 9861 1547 9919 1553
rect 9861 1513 9873 1547
rect 9907 1544 9919 1547
rect 10410 1544 10416 1556
rect 9907 1516 10416 1544
rect 9907 1513 9919 1516
rect 9861 1507 9919 1513
rect 10410 1504 10416 1516
rect 10468 1504 10474 1556
rect 10873 1547 10931 1553
rect 10873 1513 10885 1547
rect 10919 1544 10931 1547
rect 11514 1544 11520 1556
rect 10919 1516 11520 1544
rect 10919 1513 10931 1516
rect 10873 1507 10931 1513
rect 11514 1504 11520 1516
rect 11572 1504 11578 1556
rect 12345 1547 12403 1553
rect 12345 1513 12357 1547
rect 12391 1544 12403 1547
rect 12894 1544 12900 1556
rect 12391 1516 12900 1544
rect 12391 1513 12403 1516
rect 12345 1507 12403 1513
rect 12894 1504 12900 1516
rect 12952 1504 12958 1556
rect 13173 1547 13231 1553
rect 13173 1513 13185 1547
rect 13219 1544 13231 1547
rect 13630 1544 13636 1556
rect 13219 1516 13636 1544
rect 13219 1513 13231 1516
rect 13173 1507 13231 1513
rect 13630 1504 13636 1516
rect 13688 1504 13694 1556
rect 13906 1504 13912 1556
rect 13964 1504 13970 1556
rect 14461 1547 14519 1553
rect 14461 1513 14473 1547
rect 14507 1544 14519 1547
rect 14918 1544 14924 1556
rect 14507 1516 14924 1544
rect 14507 1513 14519 1516
rect 14461 1507 14519 1513
rect 14918 1504 14924 1516
rect 14976 1504 14982 1556
rect 15657 1547 15715 1553
rect 15657 1513 15669 1547
rect 15703 1544 15715 1547
rect 16114 1544 16120 1556
rect 15703 1516 16120 1544
rect 15703 1513 15715 1516
rect 15657 1507 15715 1513
rect 16114 1504 16120 1516
rect 16172 1504 16178 1556
rect 18141 1547 18199 1553
rect 18141 1513 18153 1547
rect 18187 1544 18199 1547
rect 18598 1544 18604 1556
rect 18187 1516 18604 1544
rect 18187 1513 18199 1516
rect 18141 1507 18199 1513
rect 18598 1504 18604 1516
rect 18656 1504 18662 1556
rect 20165 1547 20223 1553
rect 20165 1513 20177 1547
rect 20211 1544 20223 1547
rect 20530 1544 20536 1556
rect 20211 1516 20536 1544
rect 20211 1513 20223 1516
rect 20165 1507 20223 1513
rect 20530 1504 20536 1516
rect 20588 1504 20594 1556
rect 21821 1547 21879 1553
rect 21821 1513 21833 1547
rect 21867 1544 21879 1547
rect 22278 1544 22284 1556
rect 21867 1516 22284 1544
rect 21867 1513 21879 1516
rect 21821 1507 21879 1513
rect 22278 1504 22284 1516
rect 22336 1504 22342 1556
rect 22554 1504 22560 1556
rect 22612 1504 22618 1556
rect 22833 1547 22891 1553
rect 22833 1513 22845 1547
rect 22879 1544 22891 1547
rect 23566 1544 23572 1556
rect 22879 1516 23572 1544
rect 22879 1513 22891 1516
rect 22833 1507 22891 1513
rect 23566 1504 23572 1516
rect 23624 1504 23630 1556
rect 23753 1547 23811 1553
rect 23753 1513 23765 1547
rect 23799 1544 23811 1547
rect 24302 1544 24308 1556
rect 23799 1516 24308 1544
rect 23799 1513 23811 1516
rect 23753 1507 23811 1513
rect 24302 1504 24308 1516
rect 24360 1504 24366 1556
rect 13449 1479 13507 1485
rect 13449 1445 13461 1479
rect 13495 1476 13507 1479
rect 13924 1476 13952 1504
rect 13495 1448 13952 1476
rect 21361 1479 21419 1485
rect 13495 1445 13507 1448
rect 13449 1439 13507 1445
rect 21361 1445 21373 1479
rect 21407 1445 21419 1479
rect 21361 1439 21419 1445
rect 22097 1479 22155 1485
rect 22097 1445 22109 1479
rect 22143 1476 22155 1479
rect 22572 1476 22600 1504
rect 22143 1448 22600 1476
rect 23477 1479 23535 1485
rect 22143 1445 22155 1448
rect 22097 1439 22155 1445
rect 23477 1445 23489 1479
rect 23523 1476 23535 1479
rect 24026 1476 24032 1488
rect 23523 1448 24032 1476
rect 23523 1445 23535 1448
rect 23477 1439 23535 1445
rect 13262 1368 13268 1420
rect 13320 1408 13326 1420
rect 21376 1408 21404 1439
rect 24026 1436 24032 1448
rect 24084 1436 24090 1488
rect 13320 1380 13860 1408
rect 21376 1380 21680 1408
rect 13320 1368 13326 1380
rect 934 1300 940 1352
rect 992 1340 998 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 992 1312 1409 1340
rect 992 1300 998 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 2222 1300 2228 1352
rect 2280 1300 2286 1352
rect 3418 1300 3424 1352
rect 3476 1300 3482 1352
rect 4798 1300 4804 1352
rect 4856 1300 4862 1352
rect 5994 1300 6000 1352
rect 6052 1300 6058 1352
rect 7377 1343 7435 1349
rect 7377 1309 7389 1343
rect 7423 1340 7435 1343
rect 7423 1312 7512 1340
rect 7423 1309 7435 1312
rect 7377 1303 7435 1309
rect 3620 1244 6914 1272
rect 1578 1164 1584 1216
rect 1636 1164 1642 1216
rect 2406 1164 2412 1216
rect 2464 1164 2470 1216
rect 3620 1213 3648 1244
rect 3605 1207 3663 1213
rect 3605 1173 3617 1207
rect 3651 1173 3663 1207
rect 3605 1167 3663 1173
rect 4614 1164 4620 1216
rect 4672 1164 4678 1216
rect 5810 1164 5816 1216
rect 5868 1164 5874 1216
rect 6886 1204 6914 1244
rect 7374 1204 7380 1216
rect 6886 1176 7380 1204
rect 7374 1164 7380 1176
rect 7432 1164 7438 1216
rect 7484 1213 7512 1312
rect 7650 1300 7656 1352
rect 7708 1300 7714 1352
rect 8573 1343 8631 1349
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 8619 1312 8984 1340
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 8956 1213 8984 1312
rect 9122 1300 9128 1352
rect 9180 1300 9186 1352
rect 9769 1343 9827 1349
rect 9769 1309 9781 1343
rect 9815 1309 9827 1343
rect 9769 1303 9827 1309
rect 9784 1272 9812 1303
rect 10042 1300 10048 1352
rect 10100 1300 10106 1352
rect 10318 1300 10324 1352
rect 10376 1300 10382 1352
rect 10778 1300 10784 1352
rect 10836 1300 10842 1352
rect 11057 1343 11115 1349
rect 11057 1309 11069 1343
rect 11103 1309 11115 1343
rect 11057 1303 11115 1309
rect 11072 1272 11100 1303
rect 11974 1300 11980 1352
rect 12032 1300 12038 1352
rect 12253 1343 12311 1349
rect 12253 1309 12265 1343
rect 12299 1309 12311 1343
rect 12253 1303 12311 1309
rect 12268 1272 12296 1303
rect 12526 1300 12532 1352
rect 12584 1300 12590 1352
rect 13357 1343 13415 1349
rect 13357 1309 13369 1343
rect 13403 1309 13415 1343
rect 13357 1303 13415 1309
rect 9784 1244 10180 1272
rect 10152 1213 10180 1244
rect 10612 1244 11100 1272
rect 11808 1244 12296 1272
rect 13372 1272 13400 1303
rect 13630 1300 13636 1352
rect 13688 1300 13694 1352
rect 13832 1340 13860 1380
rect 13909 1343 13967 1349
rect 13909 1340 13921 1343
rect 13832 1312 13921 1340
rect 13909 1309 13921 1312
rect 13955 1309 13967 1343
rect 13909 1303 13967 1309
rect 14366 1300 14372 1352
rect 14424 1300 14430 1352
rect 14645 1343 14703 1349
rect 14645 1309 14657 1343
rect 14691 1309 14703 1343
rect 14645 1303 14703 1309
rect 14660 1272 14688 1303
rect 15010 1300 15016 1352
rect 15068 1300 15074 1352
rect 15378 1340 15384 1352
rect 15120 1312 15384 1340
rect 13372 1244 13768 1272
rect 10612 1213 10640 1244
rect 11808 1213 11836 1244
rect 7469 1207 7527 1213
rect 7469 1173 7481 1207
rect 7515 1173 7527 1207
rect 7469 1167 7527 1173
rect 8941 1207 8999 1213
rect 8941 1173 8953 1207
rect 8987 1173 8999 1207
rect 8941 1167 8999 1173
rect 10137 1207 10195 1213
rect 10137 1173 10149 1207
rect 10183 1173 10195 1207
rect 10137 1167 10195 1173
rect 10597 1207 10655 1213
rect 10597 1173 10609 1207
rect 10643 1173 10655 1207
rect 10597 1167 10655 1173
rect 11793 1207 11851 1213
rect 11793 1173 11805 1207
rect 11839 1173 11851 1207
rect 11793 1167 11851 1173
rect 12069 1207 12127 1213
rect 12069 1173 12081 1207
rect 12115 1204 12127 1207
rect 12618 1204 12624 1216
rect 12115 1176 12624 1204
rect 12115 1173 12127 1176
rect 12069 1167 12127 1173
rect 12618 1164 12624 1176
rect 12676 1164 12682 1216
rect 13740 1213 13768 1244
rect 14200 1244 14688 1272
rect 14200 1213 14228 1244
rect 13725 1207 13783 1213
rect 13725 1173 13737 1207
rect 13771 1173 13783 1207
rect 13725 1167 13783 1173
rect 14185 1207 14243 1213
rect 14185 1173 14197 1207
rect 14231 1173 14243 1207
rect 14185 1167 14243 1173
rect 14829 1207 14887 1213
rect 14829 1173 14841 1207
rect 14875 1204 14887 1207
rect 15120 1204 15148 1312
rect 15378 1300 15384 1312
rect 15436 1300 15442 1352
rect 15562 1300 15568 1352
rect 15620 1300 15626 1352
rect 15841 1343 15899 1349
rect 15841 1309 15853 1343
rect 15887 1309 15899 1343
rect 15841 1303 15899 1309
rect 15856 1272 15884 1303
rect 16666 1300 16672 1352
rect 16724 1300 16730 1352
rect 16942 1300 16948 1352
rect 17000 1300 17006 1352
rect 17126 1300 17132 1352
rect 17184 1300 17190 1352
rect 17954 1300 17960 1352
rect 18012 1300 18018 1352
rect 18325 1343 18383 1349
rect 18325 1309 18337 1343
rect 18371 1309 18383 1343
rect 18325 1303 18383 1309
rect 15396 1244 15884 1272
rect 15396 1213 15424 1244
rect 14875 1176 15148 1204
rect 15381 1207 15439 1213
rect 14875 1173 14887 1176
rect 14829 1167 14887 1173
rect 15381 1173 15393 1207
rect 15427 1173 15439 1207
rect 15381 1167 15439 1173
rect 16850 1164 16856 1216
rect 16908 1164 16914 1216
rect 16960 1213 16988 1300
rect 18340 1272 18368 1303
rect 19426 1300 19432 1352
rect 19484 1300 19490 1352
rect 20346 1300 20352 1352
rect 20404 1300 20410 1352
rect 21542 1300 21548 1352
rect 21600 1300 21606 1352
rect 21652 1340 21680 1380
rect 22005 1343 22063 1349
rect 22005 1340 22017 1343
rect 21652 1312 22017 1340
rect 22005 1309 22017 1312
rect 22051 1309 22063 1343
rect 22281 1343 22339 1349
rect 22281 1340 22293 1343
rect 22005 1303 22063 1309
rect 22112 1312 22293 1340
rect 17788 1244 18368 1272
rect 17788 1213 17816 1244
rect 16945 1207 17003 1213
rect 16945 1173 16957 1207
rect 16991 1173 17003 1207
rect 16945 1167 17003 1173
rect 17773 1207 17831 1213
rect 17773 1173 17785 1207
rect 17819 1173 17831 1207
rect 17773 1167 17831 1173
rect 19245 1207 19303 1213
rect 19245 1173 19257 1207
rect 19291 1204 19303 1207
rect 22112 1204 22140 1312
rect 22281 1309 22293 1312
rect 22327 1309 22339 1343
rect 22281 1303 22339 1309
rect 22738 1300 22744 1352
rect 22796 1300 22802 1352
rect 23017 1343 23075 1349
rect 23017 1309 23029 1343
rect 23063 1309 23075 1343
rect 23017 1303 23075 1309
rect 23385 1343 23443 1349
rect 23385 1309 23397 1343
rect 23431 1340 23443 1343
rect 23566 1340 23572 1352
rect 23431 1312 23572 1340
rect 23431 1309 23443 1312
rect 23385 1303 23443 1309
rect 23032 1272 23060 1303
rect 23566 1300 23572 1312
rect 23624 1300 23630 1352
rect 23661 1343 23719 1349
rect 23661 1309 23673 1343
rect 23707 1309 23719 1343
rect 23661 1303 23719 1309
rect 23937 1343 23995 1349
rect 23937 1309 23949 1343
rect 23983 1340 23995 1343
rect 23983 1312 24072 1340
rect 23983 1309 23995 1312
rect 23937 1303 23995 1309
rect 23676 1272 23704 1303
rect 22572 1244 23060 1272
rect 23216 1244 23704 1272
rect 22572 1213 22600 1244
rect 23216 1213 23244 1244
rect 24044 1213 24072 1312
rect 24210 1300 24216 1352
rect 24268 1300 24274 1352
rect 19291 1176 22140 1204
rect 22557 1207 22615 1213
rect 19291 1173 19303 1176
rect 19245 1167 19303 1173
rect 22557 1173 22569 1207
rect 22603 1173 22615 1207
rect 22557 1167 22615 1173
rect 23201 1207 23259 1213
rect 23201 1173 23213 1207
rect 23247 1173 23259 1207
rect 23201 1167 23259 1173
rect 24029 1207 24087 1213
rect 24029 1173 24041 1207
rect 24075 1173 24087 1207
rect 24029 1167 24087 1173
rect 1104 1114 25000 1136
rect 1104 1062 6884 1114
rect 6936 1062 6948 1114
rect 7000 1062 7012 1114
rect 7064 1062 7076 1114
rect 7128 1062 7140 1114
rect 7192 1062 12818 1114
rect 12870 1062 12882 1114
rect 12934 1062 12946 1114
rect 12998 1062 13010 1114
rect 13062 1062 13074 1114
rect 13126 1062 18752 1114
rect 18804 1062 18816 1114
rect 18868 1062 18880 1114
rect 18932 1062 18944 1114
rect 18996 1062 19008 1114
rect 19060 1062 24686 1114
rect 24738 1062 24750 1114
rect 24802 1062 24814 1114
rect 24866 1062 24878 1114
rect 24930 1062 24942 1114
rect 24994 1062 25000 1114
rect 1104 1040 25000 1062
rect 1578 960 1584 1012
rect 1636 960 1642 1012
rect 4614 960 4620 1012
rect 4672 1000 4678 1012
rect 7282 1000 7288 1012
rect 4672 972 7288 1000
rect 4672 960 4678 972
rect 7282 960 7288 972
rect 7340 960 7346 1012
rect 7374 960 7380 1012
rect 7432 1000 7438 1012
rect 15010 1000 15016 1012
rect 7432 972 15016 1000
rect 7432 960 7438 972
rect 15010 960 15016 972
rect 15068 960 15074 1012
rect 16666 960 16672 1012
rect 16724 960 16730 1012
rect 16850 960 16856 1012
rect 16908 1000 16914 1012
rect 20162 1000 20168 1012
rect 16908 972 20168 1000
rect 16908 960 16914 972
rect 20162 960 20168 972
rect 20220 960 20226 1012
rect 1596 932 1624 960
rect 16684 932 16712 960
rect 1596 904 16712 932
rect 2406 824 2412 876
rect 2464 824 2470 876
rect 5810 824 5816 876
rect 5868 864 5874 876
rect 10042 864 10048 876
rect 5868 836 6914 864
rect 5868 824 5874 836
rect 2424 660 2452 824
rect 6886 728 6914 836
rect 7392 836 10048 864
rect 7392 728 7420 836
rect 10042 824 10048 836
rect 10100 824 10106 876
rect 13630 864 13636 876
rect 12406 836 13636 864
rect 6886 700 7420 728
rect 8478 688 8484 740
rect 8536 728 8542 740
rect 9122 728 9128 740
rect 8536 700 9128 728
rect 8536 688 8542 700
rect 9122 688 9128 700
rect 9180 688 9186 740
rect 9674 688 9680 740
rect 9732 728 9738 740
rect 10318 728 10324 740
rect 9732 700 10324 728
rect 9732 688 9738 700
rect 10318 688 10324 700
rect 10376 688 10382 740
rect 12406 660 12434 836
rect 13630 824 13636 836
rect 13688 824 13694 876
rect 23566 688 23572 740
rect 23624 728 23630 740
rect 24854 728 24860 740
rect 23624 700 24860 728
rect 23624 688 23630 700
rect 24854 688 24860 700
rect 24912 688 24918 740
rect 2424 632 12434 660
rect 7282 552 7288 604
rect 7340 592 7346 604
rect 12526 592 12532 604
rect 7340 564 12532 592
rect 7340 552 7346 564
rect 12526 552 12532 564
rect 12584 552 12590 604
<< via1 >>
rect 7840 9936 7892 9988
rect 18604 9936 18656 9988
rect 18512 9868 18564 9920
rect 15016 9800 15068 9852
rect 6644 9732 6696 9784
rect 7472 9732 7524 9784
rect 10600 9732 10652 9784
rect 14096 9732 14148 9784
rect 3700 9664 3752 9716
rect 15200 9664 15252 9716
rect 7564 9596 7616 9648
rect 18236 9596 18288 9648
rect 2872 9528 2924 9580
rect 11612 9528 11664 9580
rect 11704 9528 11756 9580
rect 19984 9528 20036 9580
rect 8944 9460 8996 9512
rect 16304 9460 16356 9512
rect 8392 9392 8444 9444
rect 13544 9392 13596 9444
rect 2504 9324 2556 9376
rect 11428 9324 11480 9376
rect 11612 9324 11664 9376
rect 14188 9324 14240 9376
rect 2780 9256 2832 9308
rect 13912 9256 13964 9308
rect 2320 9188 2372 9240
rect 1768 9120 1820 9172
rect 3700 9120 3752 9172
rect 8024 9188 8076 9240
rect 17500 9188 17552 9240
rect 12624 9120 12676 9172
rect 18696 9120 18748 9172
rect 19708 9120 19760 9172
rect 9404 9052 9456 9104
rect 16672 9052 16724 9104
rect 21732 9052 21784 9104
rect 22928 9052 22980 9104
rect 5540 8848 5592 8900
rect 8668 8848 8720 8900
rect 16948 8984 17000 9036
rect 17224 8916 17276 8968
rect 15844 8848 15896 8900
rect 3148 8780 3200 8832
rect 8392 8780 8444 8832
rect 9220 8780 9272 8832
rect 9956 8780 10008 8832
rect 11152 8780 11204 8832
rect 12716 8780 12768 8832
rect 14740 8780 14792 8832
rect 6884 8678 6936 8730
rect 6948 8678 7000 8730
rect 7012 8678 7064 8730
rect 7076 8678 7128 8730
rect 7140 8678 7192 8730
rect 12818 8678 12870 8730
rect 12882 8678 12934 8730
rect 12946 8678 12998 8730
rect 13010 8678 13062 8730
rect 13074 8678 13126 8730
rect 18752 8678 18804 8730
rect 18816 8678 18868 8730
rect 18880 8678 18932 8730
rect 18944 8678 18996 8730
rect 19008 8678 19060 8730
rect 24686 8678 24738 8730
rect 24750 8678 24802 8730
rect 24814 8678 24866 8730
rect 24878 8678 24930 8730
rect 24942 8678 24994 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 2964 8576 3016 8628
rect 664 8508 716 8560
rect 4344 8576 4396 8628
rect 5172 8576 5224 8628
rect 5448 8576 5500 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 6736 8576 6788 8628
rect 7656 8576 7708 8628
rect 8116 8576 8168 8628
rect 8484 8576 8536 8628
rect 8760 8576 8812 8628
rect 9036 8576 9088 8628
rect 9312 8576 9364 8628
rect 11428 8576 11480 8628
rect 12164 8576 12216 8628
rect 12624 8576 12676 8628
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 14188 8576 14240 8628
rect 14464 8576 14516 8628
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 2780 8440 2832 8492
rect 7840 8508 7892 8560
rect 8024 8551 8076 8560
rect 8024 8517 8033 8551
rect 8033 8517 8067 8551
rect 8067 8517 8076 8551
rect 8024 8508 8076 8517
rect 5540 8440 5592 8492
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 6644 8440 6696 8492
rect 7472 8440 7524 8492
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 8392 8440 8444 8492
rect 9956 8508 10008 8560
rect 9220 8440 9272 8492
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 10600 8440 10652 8492
rect 11152 8440 11204 8492
rect 11520 8440 11572 8492
rect 7472 8304 7524 8356
rect 7564 8304 7616 8356
rect 9772 8372 9824 8424
rect 9864 8372 9916 8424
rect 9588 8304 9640 8356
rect 5908 8236 5960 8288
rect 8392 8236 8444 8288
rect 8484 8236 8536 8288
rect 9956 8236 10008 8288
rect 11060 8304 11112 8356
rect 11336 8236 11388 8288
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 12532 8487 12584 8492
rect 12532 8453 12541 8487
rect 12541 8453 12575 8487
rect 12575 8453 12584 8487
rect 12532 8440 12584 8453
rect 12716 8440 12768 8492
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 13544 8440 13596 8492
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 13636 8440 13688 8449
rect 12440 8372 12492 8424
rect 12808 8372 12860 8424
rect 14004 8508 14056 8560
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 14464 8440 14516 8492
rect 15200 8619 15252 8628
rect 15200 8585 15209 8619
rect 15209 8585 15243 8619
rect 15243 8585 15252 8619
rect 15200 8576 15252 8585
rect 15476 8576 15528 8628
rect 15844 8619 15896 8628
rect 15844 8585 15853 8619
rect 15853 8585 15887 8619
rect 15887 8585 15896 8619
rect 15844 8576 15896 8585
rect 16304 8576 16356 8628
rect 16396 8576 16448 8628
rect 16672 8619 16724 8628
rect 16672 8585 16681 8619
rect 16681 8585 16715 8619
rect 16715 8585 16724 8619
rect 16672 8576 16724 8585
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 17224 8619 17276 8628
rect 17224 8585 17233 8619
rect 17233 8585 17267 8619
rect 17267 8585 17276 8619
rect 17224 8576 17276 8585
rect 17500 8619 17552 8628
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 17592 8576 17644 8628
rect 15200 8440 15252 8492
rect 14556 8372 14608 8424
rect 15660 8440 15712 8492
rect 14372 8304 14424 8356
rect 14464 8347 14516 8356
rect 14464 8313 14473 8347
rect 14473 8313 14507 8347
rect 14507 8313 14516 8347
rect 14464 8304 14516 8313
rect 15384 8304 15436 8356
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 16672 8372 16724 8424
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17224 8372 17276 8424
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 18604 8576 18656 8628
rect 19984 8619 20036 8628
rect 19984 8585 19993 8619
rect 19993 8585 20027 8619
rect 20027 8585 20036 8619
rect 19984 8576 20036 8585
rect 20076 8576 20128 8628
rect 20536 8576 20588 8628
rect 20904 8576 20956 8628
rect 21548 8576 21600 8628
rect 22928 8619 22980 8628
rect 22928 8585 22937 8619
rect 22937 8585 22971 8619
rect 22971 8585 22980 8619
rect 22928 8576 22980 8585
rect 23112 8576 23164 8628
rect 18972 8508 19024 8560
rect 19156 8508 19208 8560
rect 14556 8236 14608 8288
rect 14740 8279 14792 8288
rect 14740 8245 14749 8279
rect 14749 8245 14783 8279
rect 14783 8245 14792 8279
rect 14740 8236 14792 8245
rect 15016 8236 15068 8288
rect 17868 8236 17920 8288
rect 18236 8347 18288 8356
rect 18236 8313 18245 8347
rect 18245 8313 18279 8347
rect 18279 8313 18288 8347
rect 18236 8304 18288 8313
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 18604 8372 18656 8424
rect 19708 8483 19760 8492
rect 19708 8449 19717 8483
rect 19717 8449 19751 8483
rect 19751 8449 19760 8483
rect 19708 8440 19760 8449
rect 20168 8483 20220 8492
rect 20168 8449 20177 8483
rect 20177 8449 20211 8483
rect 20211 8449 20220 8483
rect 20168 8440 20220 8449
rect 20812 8440 20864 8492
rect 21272 8440 21324 8492
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 22468 8440 22520 8492
rect 22928 8440 22980 8492
rect 20996 8372 21048 8424
rect 18604 8279 18656 8288
rect 18604 8245 18613 8279
rect 18613 8245 18647 8279
rect 18647 8245 18656 8279
rect 18604 8236 18656 8245
rect 19156 8236 19208 8288
rect 19340 8236 19392 8288
rect 3917 8134 3969 8186
rect 3981 8134 4033 8186
rect 4045 8134 4097 8186
rect 4109 8134 4161 8186
rect 4173 8134 4225 8186
rect 9851 8134 9903 8186
rect 9915 8134 9967 8186
rect 9979 8134 10031 8186
rect 10043 8134 10095 8186
rect 10107 8134 10159 8186
rect 15785 8134 15837 8186
rect 15849 8134 15901 8186
rect 15913 8134 15965 8186
rect 15977 8134 16029 8186
rect 16041 8134 16093 8186
rect 21719 8134 21771 8186
rect 21783 8134 21835 8186
rect 21847 8134 21899 8186
rect 21911 8134 21963 8186
rect 21975 8134 22027 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 2412 8075 2464 8084
rect 2412 8041 2421 8075
rect 2421 8041 2455 8075
rect 2455 8041 2464 8075
rect 2412 8032 2464 8041
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 3332 8075 3384 8084
rect 3332 8041 3341 8075
rect 3341 8041 3375 8075
rect 3375 8041 3384 8075
rect 3332 8032 3384 8041
rect 4160 8075 4212 8084
rect 4160 8041 4169 8075
rect 4169 8041 4203 8075
rect 4203 8041 4212 8075
rect 4160 8032 4212 8041
rect 4988 8075 5040 8084
rect 4988 8041 4997 8075
rect 4997 8041 5031 8075
rect 5031 8041 5040 8075
rect 4988 8032 5040 8041
rect 1768 7828 1820 7880
rect 2320 7828 2372 7880
rect 3148 7828 3200 7880
rect 5908 8032 5960 8084
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 6276 8032 6328 8084
rect 6644 8075 6696 8084
rect 6644 8041 6653 8075
rect 6653 8041 6687 8075
rect 6687 8041 6696 8075
rect 6644 8032 6696 8041
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 7380 8032 7432 8084
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 8392 8032 8444 8084
rect 11152 8032 11204 8084
rect 5356 7896 5408 7948
rect 9680 7964 9732 8016
rect 5816 7828 5868 7880
rect 7932 7896 7984 7948
rect 8576 7896 8628 7948
rect 8944 7828 8996 7880
rect 3240 7692 3292 7744
rect 5448 7760 5500 7812
rect 6552 7803 6604 7812
rect 6552 7769 6561 7803
rect 6561 7769 6595 7803
rect 6595 7769 6604 7803
rect 6552 7760 6604 7769
rect 8116 7760 8168 7812
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 9772 7828 9824 7880
rect 10876 7964 10928 8016
rect 10600 7896 10652 7948
rect 11520 7964 11572 8016
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 12164 7896 12216 7948
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 12992 8075 13044 8084
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 14096 8032 14148 8084
rect 14188 8032 14240 8084
rect 15200 8075 15252 8084
rect 15200 8041 15209 8075
rect 15209 8041 15243 8075
rect 15243 8041 15252 8075
rect 15200 8032 15252 8041
rect 15660 8032 15712 8084
rect 16856 8032 16908 8084
rect 17408 8032 17460 8084
rect 17776 8032 17828 8084
rect 17868 8032 17920 8084
rect 16488 7964 16540 8016
rect 12348 7828 12400 7880
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 14832 7828 14884 7880
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 16212 7896 16264 7948
rect 15660 7760 15712 7812
rect 16120 7828 16172 7880
rect 17224 8007 17276 8016
rect 17224 7973 17233 8007
rect 17233 7973 17267 8007
rect 17267 7973 17276 8007
rect 17224 7964 17276 7973
rect 17316 7964 17368 8016
rect 17040 7896 17092 7948
rect 18604 8032 18656 8084
rect 18880 8032 18932 8084
rect 19340 8032 19392 8084
rect 21180 8032 21232 8084
rect 22560 8075 22612 8084
rect 22560 8041 22569 8075
rect 22569 8041 22603 8075
rect 22603 8041 22612 8075
rect 22560 8032 22612 8041
rect 22836 8032 22888 8084
rect 23388 8032 23440 8084
rect 23664 8032 23716 8084
rect 18788 7964 18840 8016
rect 16764 7760 16816 7812
rect 18144 7828 18196 7880
rect 19156 7828 19208 7880
rect 19340 7871 19392 7880
rect 19340 7837 19349 7871
rect 19349 7837 19383 7871
rect 19383 7837 19392 7871
rect 19340 7828 19392 7837
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 25596 7828 25648 7880
rect 10048 7692 10100 7744
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 10784 7735 10836 7744
rect 10784 7701 10793 7735
rect 10793 7701 10827 7735
rect 10827 7701 10836 7735
rect 10784 7692 10836 7701
rect 10876 7692 10928 7744
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 18052 7692 18104 7744
rect 19524 7735 19576 7744
rect 19524 7701 19533 7735
rect 19533 7701 19567 7735
rect 19567 7701 19576 7735
rect 19524 7692 19576 7701
rect 19800 7735 19852 7744
rect 19800 7701 19809 7735
rect 19809 7701 19843 7735
rect 19843 7701 19852 7735
rect 19800 7692 19852 7701
rect 20076 7735 20128 7744
rect 20076 7701 20085 7735
rect 20085 7701 20119 7735
rect 20119 7701 20128 7735
rect 20076 7692 20128 7701
rect 21916 7803 21968 7812
rect 21916 7769 21925 7803
rect 21925 7769 21959 7803
rect 21959 7769 21968 7803
rect 21916 7760 21968 7769
rect 22468 7803 22520 7812
rect 22468 7769 22477 7803
rect 22477 7769 22511 7803
rect 22511 7769 22520 7803
rect 22468 7760 22520 7769
rect 22652 7760 22704 7812
rect 23848 7803 23900 7812
rect 23848 7769 23857 7803
rect 23857 7769 23891 7803
rect 23891 7769 23900 7803
rect 23848 7760 23900 7769
rect 23756 7692 23808 7744
rect 6884 7590 6936 7642
rect 6948 7590 7000 7642
rect 7012 7590 7064 7642
rect 7076 7590 7128 7642
rect 7140 7590 7192 7642
rect 12818 7590 12870 7642
rect 12882 7590 12934 7642
rect 12946 7590 12998 7642
rect 13010 7590 13062 7642
rect 13074 7590 13126 7642
rect 18752 7590 18804 7642
rect 18816 7590 18868 7642
rect 18880 7590 18932 7642
rect 18944 7590 18996 7642
rect 19008 7590 19060 7642
rect 24686 7590 24738 7642
rect 24750 7590 24802 7642
rect 24814 7590 24866 7642
rect 24878 7590 24930 7642
rect 24942 7590 24994 7642
rect 1308 7488 1360 7540
rect 2228 7488 2280 7540
rect 3792 7488 3844 7540
rect 4620 7531 4672 7540
rect 4620 7497 4629 7531
rect 4629 7497 4663 7531
rect 4663 7497 4672 7531
rect 4620 7488 4672 7497
rect 5356 7488 5408 7540
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 5632 7488 5684 7540
rect 5816 7488 5868 7540
rect 6552 7488 6604 7540
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 7840 7488 7892 7540
rect 8668 7488 8720 7540
rect 9680 7488 9732 7540
rect 10324 7488 10376 7540
rect 11152 7488 11204 7540
rect 17776 7488 17828 7540
rect 21916 7488 21968 7540
rect 22560 7488 22612 7540
rect 24216 7488 24268 7540
rect 25320 7488 25372 7540
rect 1952 7463 2004 7472
rect 1952 7429 1961 7463
rect 1961 7429 1995 7463
rect 1995 7429 2004 7463
rect 1952 7420 2004 7429
rect 2688 7420 2740 7472
rect 3516 7148 3568 7200
rect 19800 7420 19852 7472
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 7564 7352 7616 7404
rect 7380 7284 7432 7336
rect 8668 7352 8720 7404
rect 10324 7352 10376 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 10784 7352 10836 7404
rect 20720 7352 20772 7404
rect 23112 7395 23164 7404
rect 23112 7361 23121 7395
rect 23121 7361 23155 7395
rect 23155 7361 23164 7395
rect 23112 7352 23164 7361
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 23664 7352 23716 7361
rect 23296 7284 23348 7336
rect 25044 7284 25096 7336
rect 6276 7148 6328 7200
rect 6368 7191 6420 7200
rect 6368 7157 6377 7191
rect 6377 7157 6411 7191
rect 6411 7157 6420 7191
rect 6368 7148 6420 7157
rect 10508 7216 10560 7268
rect 10600 7216 10652 7268
rect 8484 7148 8536 7200
rect 8668 7148 8720 7200
rect 3917 7046 3969 7098
rect 3981 7046 4033 7098
rect 4045 7046 4097 7098
rect 4109 7046 4161 7098
rect 4173 7046 4225 7098
rect 9851 7046 9903 7098
rect 9915 7046 9967 7098
rect 9979 7046 10031 7098
rect 10043 7046 10095 7098
rect 10107 7046 10159 7098
rect 15785 7046 15837 7098
rect 15849 7046 15901 7098
rect 15913 7046 15965 7098
rect 15977 7046 16029 7098
rect 16041 7046 16093 7098
rect 21719 7046 21771 7098
rect 21783 7046 21835 7098
rect 21847 7046 21899 7098
rect 21911 7046 21963 7098
rect 21975 7046 22027 7098
rect 3240 6944 3292 6996
rect 11060 6944 11112 6996
rect 11336 6944 11388 6996
rect 6276 6876 6328 6928
rect 1032 6808 1084 6860
rect 8116 6808 8168 6860
rect 18052 6944 18104 6996
rect 22100 6944 22152 6996
rect 24584 6808 24636 6860
rect 9772 6740 9824 6792
rect 22100 6740 22152 6792
rect 7748 6672 7800 6724
rect 23020 6715 23072 6724
rect 23020 6681 23029 6715
rect 23029 6681 23063 6715
rect 23063 6681 23072 6715
rect 23020 6672 23072 6681
rect 204 6604 256 6656
rect 6884 6502 6936 6554
rect 6948 6502 7000 6554
rect 7012 6502 7064 6554
rect 7076 6502 7128 6554
rect 7140 6502 7192 6554
rect 12818 6502 12870 6554
rect 12882 6502 12934 6554
rect 12946 6502 12998 6554
rect 13010 6502 13062 6554
rect 13074 6502 13126 6554
rect 18752 6502 18804 6554
rect 18816 6502 18868 6554
rect 18880 6502 18932 6554
rect 18944 6502 18996 6554
rect 19008 6502 19060 6554
rect 24686 6502 24738 6554
rect 24750 6502 24802 6554
rect 24814 6502 24866 6554
rect 24878 6502 24930 6554
rect 24942 6502 24994 6554
rect 756 6400 808 6452
rect 23940 6400 23992 6452
rect 24492 6400 24544 6452
rect 6368 6332 6420 6384
rect 23388 6332 23440 6384
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 23480 6307 23532 6316
rect 23480 6273 23489 6307
rect 23489 6273 23523 6307
rect 23523 6273 23532 6307
rect 23480 6264 23532 6273
rect 23848 6060 23900 6112
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 9851 5958 9903 6010
rect 9915 5958 9967 6010
rect 9979 5958 10031 6010
rect 10043 5958 10095 6010
rect 10107 5958 10159 6010
rect 15785 5958 15837 6010
rect 15849 5958 15901 6010
rect 15913 5958 15965 6010
rect 15977 5958 16029 6010
rect 16041 5958 16093 6010
rect 21719 5958 21771 6010
rect 21783 5958 21835 6010
rect 21847 5958 21899 6010
rect 21911 5958 21963 6010
rect 21975 5958 22027 6010
rect 17500 5856 17552 5908
rect 16948 5695 17000 5704
rect 16948 5661 16957 5695
rect 16957 5661 16991 5695
rect 16991 5661 17000 5695
rect 16948 5652 17000 5661
rect 6884 5414 6936 5466
rect 6948 5414 7000 5466
rect 7012 5414 7064 5466
rect 7076 5414 7128 5466
rect 7140 5414 7192 5466
rect 12818 5414 12870 5466
rect 12882 5414 12934 5466
rect 12946 5414 12998 5466
rect 13010 5414 13062 5466
rect 13074 5414 13126 5466
rect 18752 5414 18804 5466
rect 18816 5414 18868 5466
rect 18880 5414 18932 5466
rect 18944 5414 18996 5466
rect 19008 5414 19060 5466
rect 24686 5414 24738 5466
rect 24750 5414 24802 5466
rect 24814 5414 24866 5466
rect 24878 5414 24930 5466
rect 24942 5414 24994 5466
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 9851 4870 9903 4922
rect 9915 4870 9967 4922
rect 9979 4870 10031 4922
rect 10043 4870 10095 4922
rect 10107 4870 10159 4922
rect 15785 4870 15837 4922
rect 15849 4870 15901 4922
rect 15913 4870 15965 4922
rect 15977 4870 16029 4922
rect 16041 4870 16093 4922
rect 21719 4870 21771 4922
rect 21783 4870 21835 4922
rect 21847 4870 21899 4922
rect 21911 4870 21963 4922
rect 21975 4870 22027 4922
rect 6884 4326 6936 4378
rect 6948 4326 7000 4378
rect 7012 4326 7064 4378
rect 7076 4326 7128 4378
rect 7140 4326 7192 4378
rect 12818 4326 12870 4378
rect 12882 4326 12934 4378
rect 12946 4326 12998 4378
rect 13010 4326 13062 4378
rect 13074 4326 13126 4378
rect 18752 4326 18804 4378
rect 18816 4326 18868 4378
rect 18880 4326 18932 4378
rect 18944 4326 18996 4378
rect 19008 4326 19060 4378
rect 24686 4326 24738 4378
rect 24750 4326 24802 4378
rect 24814 4326 24866 4378
rect 24878 4326 24930 4378
rect 24942 4326 24994 4378
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 9851 3782 9903 3834
rect 9915 3782 9967 3834
rect 9979 3782 10031 3834
rect 10043 3782 10095 3834
rect 10107 3782 10159 3834
rect 15785 3782 15837 3834
rect 15849 3782 15901 3834
rect 15913 3782 15965 3834
rect 15977 3782 16029 3834
rect 16041 3782 16093 3834
rect 21719 3782 21771 3834
rect 21783 3782 21835 3834
rect 21847 3782 21899 3834
rect 21911 3782 21963 3834
rect 21975 3782 22027 3834
rect 6884 3238 6936 3290
rect 6948 3238 7000 3290
rect 7012 3238 7064 3290
rect 7076 3238 7128 3290
rect 7140 3238 7192 3290
rect 12818 3238 12870 3290
rect 12882 3238 12934 3290
rect 12946 3238 12998 3290
rect 13010 3238 13062 3290
rect 13074 3238 13126 3290
rect 18752 3238 18804 3290
rect 18816 3238 18868 3290
rect 18880 3238 18932 3290
rect 18944 3238 18996 3290
rect 19008 3238 19060 3290
rect 24686 3238 24738 3290
rect 24750 3238 24802 3290
rect 24814 3238 24866 3290
rect 24878 3238 24930 3290
rect 24942 3238 24994 3290
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 9851 2694 9903 2746
rect 9915 2694 9967 2746
rect 9979 2694 10031 2746
rect 10043 2694 10095 2746
rect 10107 2694 10159 2746
rect 15785 2694 15837 2746
rect 15849 2694 15901 2746
rect 15913 2694 15965 2746
rect 15977 2694 16029 2746
rect 16041 2694 16093 2746
rect 21719 2694 21771 2746
rect 21783 2694 21835 2746
rect 21847 2694 21899 2746
rect 21911 2694 21963 2746
rect 21975 2694 22027 2746
rect 13820 2592 13872 2644
rect 22652 2592 22704 2644
rect 22928 2592 22980 2644
rect 15108 2524 15160 2576
rect 13728 2388 13780 2440
rect 21272 2388 21324 2440
rect 22376 2388 22428 2440
rect 23664 2388 23716 2440
rect 23296 2320 23348 2372
rect 24124 2320 24176 2372
rect 10600 2252 10652 2304
rect 20904 2252 20956 2304
rect 6884 2150 6936 2202
rect 6948 2150 7000 2202
rect 7012 2150 7064 2202
rect 7076 2150 7128 2202
rect 7140 2150 7192 2202
rect 12818 2150 12870 2202
rect 12882 2150 12934 2202
rect 12946 2150 12998 2202
rect 13010 2150 13062 2202
rect 13074 2150 13126 2202
rect 18752 2150 18804 2202
rect 18816 2150 18868 2202
rect 18880 2150 18932 2202
rect 18944 2150 18996 2202
rect 19008 2150 19060 2202
rect 24686 2150 24738 2202
rect 24750 2150 24802 2202
rect 24814 2150 24866 2202
rect 24878 2150 24930 2202
rect 24942 2150 24994 2202
rect 9128 2091 9180 2100
rect 9128 2057 9137 2091
rect 9137 2057 9171 2091
rect 9171 2057 9180 2091
rect 9128 2048 9180 2057
rect 10232 2091 10284 2100
rect 10232 2057 10241 2091
rect 10241 2057 10275 2091
rect 10275 2057 10284 2091
rect 10232 2048 10284 2057
rect 10600 2091 10652 2100
rect 10600 2057 10609 2091
rect 10609 2057 10643 2091
rect 10643 2057 10652 2091
rect 10600 2048 10652 2057
rect 11704 2091 11756 2100
rect 11704 2057 11713 2091
rect 11713 2057 11747 2091
rect 11747 2057 11756 2091
rect 11704 2048 11756 2057
rect 13728 2048 13780 2100
rect 13820 2091 13872 2100
rect 13820 2057 13829 2091
rect 13829 2057 13863 2091
rect 13863 2057 13872 2091
rect 13820 2048 13872 2057
rect 15108 2091 15160 2100
rect 15108 2057 15117 2091
rect 15117 2057 15151 2091
rect 15151 2057 15160 2091
rect 15108 2048 15160 2057
rect 17776 2048 17828 2100
rect 22100 2091 22152 2100
rect 22100 2057 22109 2091
rect 22109 2057 22143 2091
rect 22143 2057 22152 2091
rect 22100 2048 22152 2057
rect 22376 2091 22428 2100
rect 22376 2057 22385 2091
rect 22385 2057 22419 2091
rect 22419 2057 22428 2091
rect 22376 2048 22428 2057
rect 23112 2048 23164 2100
rect 23756 2048 23808 2100
rect 24124 2091 24176 2100
rect 24124 2057 24133 2091
rect 24133 2057 24167 2091
rect 24167 2057 24176 2091
rect 24124 2048 24176 2057
rect 7748 1955 7800 1964
rect 7748 1921 7757 1955
rect 7757 1921 7791 1955
rect 7791 1921 7800 1955
rect 7748 1912 7800 1921
rect 8944 1955 8996 1964
rect 8944 1921 8953 1955
rect 8953 1921 8987 1955
rect 8987 1921 8996 1955
rect 8944 1912 8996 1921
rect 9772 1912 9824 1964
rect 10416 1955 10468 1964
rect 10416 1921 10425 1955
rect 10425 1921 10459 1955
rect 10459 1921 10468 1955
rect 10416 1912 10468 1921
rect 11520 1955 11572 1964
rect 11520 1921 11529 1955
rect 11529 1921 11563 1955
rect 11563 1921 11572 1955
rect 11520 1912 11572 1921
rect 12624 1955 12676 1964
rect 12624 1921 12633 1955
rect 12633 1921 12667 1955
rect 12667 1921 12676 1955
rect 12624 1912 12676 1921
rect 12900 1955 12952 1964
rect 12900 1921 12909 1955
rect 12909 1921 12943 1955
rect 12943 1921 12952 1955
rect 12900 1912 12952 1921
rect 13636 1955 13688 1964
rect 13636 1921 13645 1955
rect 13645 1921 13679 1955
rect 13679 1921 13688 1955
rect 13636 1912 13688 1921
rect 13912 1955 13964 1964
rect 13912 1921 13921 1955
rect 13921 1921 13955 1955
rect 13955 1921 13964 1955
rect 13912 1912 13964 1921
rect 14924 1955 14976 1964
rect 14924 1921 14933 1955
rect 14933 1921 14967 1955
rect 14967 1921 14976 1955
rect 14924 1912 14976 1921
rect 15384 1955 15436 1964
rect 15384 1921 15393 1955
rect 15393 1921 15427 1955
rect 15427 1921 15436 1955
rect 15384 1912 15436 1921
rect 16120 1955 16172 1964
rect 16120 1921 16129 1955
rect 16129 1921 16163 1955
rect 16163 1921 16172 1955
rect 16120 1912 16172 1921
rect 16304 1912 16356 1964
rect 7932 1819 7984 1828
rect 7932 1785 7941 1819
rect 7941 1785 7975 1819
rect 7975 1785 7984 1819
rect 7932 1776 7984 1785
rect 18604 1955 18656 1964
rect 18604 1921 18613 1955
rect 18613 1921 18647 1955
rect 18647 1921 18656 1955
rect 18604 1912 18656 1921
rect 20536 1955 20588 1964
rect 20536 1921 20545 1955
rect 20545 1921 20579 1955
rect 20579 1921 20588 1955
rect 20536 1912 20588 1921
rect 20720 1912 20772 1964
rect 22284 1955 22336 1964
rect 22284 1921 22293 1955
rect 22293 1921 22327 1955
rect 22327 1921 22336 1955
rect 22284 1912 22336 1921
rect 22560 1955 22612 1964
rect 22560 1921 22569 1955
rect 22569 1921 22603 1955
rect 22603 1921 22612 1955
rect 22560 1912 22612 1921
rect 23572 1912 23624 1964
rect 24032 1955 24084 1964
rect 24032 1921 24041 1955
rect 24041 1921 24075 1955
rect 24075 1921 24084 1955
rect 24032 1912 24084 1921
rect 24308 1955 24360 1964
rect 24308 1921 24317 1955
rect 24317 1921 24351 1955
rect 24351 1921 24360 1955
rect 24308 1912 24360 1921
rect 23388 1776 23440 1828
rect 23480 1776 23532 1828
rect 20812 1708 20864 1760
rect 3917 1606 3969 1658
rect 3981 1606 4033 1658
rect 4045 1606 4097 1658
rect 4109 1606 4161 1658
rect 4173 1606 4225 1658
rect 9851 1606 9903 1658
rect 9915 1606 9967 1658
rect 9979 1606 10031 1658
rect 10043 1606 10095 1658
rect 10107 1606 10159 1658
rect 15785 1606 15837 1658
rect 15849 1606 15901 1658
rect 15913 1606 15965 1658
rect 15977 1606 16029 1658
rect 16041 1606 16093 1658
rect 21719 1606 21771 1658
rect 21783 1606 21835 1658
rect 21847 1606 21899 1658
rect 21911 1606 21963 1658
rect 21975 1606 22027 1658
rect 7748 1504 7800 1556
rect 8944 1504 8996 1556
rect 9772 1504 9824 1556
rect 10416 1504 10468 1556
rect 11520 1504 11572 1556
rect 12900 1504 12952 1556
rect 13636 1504 13688 1556
rect 13912 1504 13964 1556
rect 14924 1504 14976 1556
rect 16120 1504 16172 1556
rect 18604 1504 18656 1556
rect 20536 1504 20588 1556
rect 22284 1504 22336 1556
rect 22560 1504 22612 1556
rect 23572 1504 23624 1556
rect 24308 1504 24360 1556
rect 13268 1368 13320 1420
rect 24032 1436 24084 1488
rect 940 1300 992 1352
rect 2228 1343 2280 1352
rect 2228 1309 2237 1343
rect 2237 1309 2271 1343
rect 2271 1309 2280 1343
rect 2228 1300 2280 1309
rect 3424 1343 3476 1352
rect 3424 1309 3433 1343
rect 3433 1309 3467 1343
rect 3467 1309 3476 1343
rect 3424 1300 3476 1309
rect 4804 1343 4856 1352
rect 4804 1309 4813 1343
rect 4813 1309 4847 1343
rect 4847 1309 4856 1343
rect 4804 1300 4856 1309
rect 6000 1343 6052 1352
rect 6000 1309 6009 1343
rect 6009 1309 6043 1343
rect 6043 1309 6052 1343
rect 6000 1300 6052 1309
rect 1584 1207 1636 1216
rect 1584 1173 1593 1207
rect 1593 1173 1627 1207
rect 1627 1173 1636 1207
rect 1584 1164 1636 1173
rect 2412 1207 2464 1216
rect 2412 1173 2421 1207
rect 2421 1173 2455 1207
rect 2455 1173 2464 1207
rect 2412 1164 2464 1173
rect 4620 1207 4672 1216
rect 4620 1173 4629 1207
rect 4629 1173 4663 1207
rect 4663 1173 4672 1207
rect 4620 1164 4672 1173
rect 5816 1207 5868 1216
rect 5816 1173 5825 1207
rect 5825 1173 5859 1207
rect 5859 1173 5868 1207
rect 5816 1164 5868 1173
rect 7380 1164 7432 1216
rect 7656 1343 7708 1352
rect 7656 1309 7665 1343
rect 7665 1309 7699 1343
rect 7699 1309 7708 1343
rect 7656 1300 7708 1309
rect 9128 1343 9180 1352
rect 9128 1309 9137 1343
rect 9137 1309 9171 1343
rect 9171 1309 9180 1343
rect 9128 1300 9180 1309
rect 10048 1343 10100 1352
rect 10048 1309 10057 1343
rect 10057 1309 10091 1343
rect 10091 1309 10100 1343
rect 10048 1300 10100 1309
rect 10324 1343 10376 1352
rect 10324 1309 10333 1343
rect 10333 1309 10367 1343
rect 10367 1309 10376 1343
rect 10324 1300 10376 1309
rect 10784 1343 10836 1352
rect 10784 1309 10793 1343
rect 10793 1309 10827 1343
rect 10827 1309 10836 1343
rect 10784 1300 10836 1309
rect 11980 1343 12032 1352
rect 11980 1309 11989 1343
rect 11989 1309 12023 1343
rect 12023 1309 12032 1343
rect 11980 1300 12032 1309
rect 12532 1343 12584 1352
rect 12532 1309 12541 1343
rect 12541 1309 12575 1343
rect 12575 1309 12584 1343
rect 12532 1300 12584 1309
rect 13636 1343 13688 1352
rect 13636 1309 13645 1343
rect 13645 1309 13679 1343
rect 13679 1309 13688 1343
rect 13636 1300 13688 1309
rect 14372 1343 14424 1352
rect 14372 1309 14381 1343
rect 14381 1309 14415 1343
rect 14415 1309 14424 1343
rect 14372 1300 14424 1309
rect 15016 1343 15068 1352
rect 15016 1309 15025 1343
rect 15025 1309 15059 1343
rect 15059 1309 15068 1343
rect 15016 1300 15068 1309
rect 12624 1164 12676 1216
rect 15384 1300 15436 1352
rect 15568 1343 15620 1352
rect 15568 1309 15577 1343
rect 15577 1309 15611 1343
rect 15611 1309 15620 1343
rect 15568 1300 15620 1309
rect 16672 1343 16724 1352
rect 16672 1309 16681 1343
rect 16681 1309 16715 1343
rect 16715 1309 16724 1343
rect 16672 1300 16724 1309
rect 16948 1300 17000 1352
rect 17132 1343 17184 1352
rect 17132 1309 17141 1343
rect 17141 1309 17175 1343
rect 17175 1309 17184 1343
rect 17132 1300 17184 1309
rect 17960 1343 18012 1352
rect 17960 1309 17969 1343
rect 17969 1309 18003 1343
rect 18003 1309 18012 1343
rect 17960 1300 18012 1309
rect 16856 1207 16908 1216
rect 16856 1173 16865 1207
rect 16865 1173 16899 1207
rect 16899 1173 16908 1207
rect 16856 1164 16908 1173
rect 19432 1343 19484 1352
rect 19432 1309 19441 1343
rect 19441 1309 19475 1343
rect 19475 1309 19484 1343
rect 19432 1300 19484 1309
rect 20352 1343 20404 1352
rect 20352 1309 20361 1343
rect 20361 1309 20395 1343
rect 20395 1309 20404 1343
rect 20352 1300 20404 1309
rect 21548 1343 21600 1352
rect 21548 1309 21557 1343
rect 21557 1309 21591 1343
rect 21591 1309 21600 1343
rect 21548 1300 21600 1309
rect 22744 1343 22796 1352
rect 22744 1309 22753 1343
rect 22753 1309 22787 1343
rect 22787 1309 22796 1343
rect 22744 1300 22796 1309
rect 23572 1300 23624 1352
rect 24216 1343 24268 1352
rect 24216 1309 24225 1343
rect 24225 1309 24259 1343
rect 24259 1309 24268 1343
rect 24216 1300 24268 1309
rect 6884 1062 6936 1114
rect 6948 1062 7000 1114
rect 7012 1062 7064 1114
rect 7076 1062 7128 1114
rect 7140 1062 7192 1114
rect 12818 1062 12870 1114
rect 12882 1062 12934 1114
rect 12946 1062 12998 1114
rect 13010 1062 13062 1114
rect 13074 1062 13126 1114
rect 18752 1062 18804 1114
rect 18816 1062 18868 1114
rect 18880 1062 18932 1114
rect 18944 1062 18996 1114
rect 19008 1062 19060 1114
rect 24686 1062 24738 1114
rect 24750 1062 24802 1114
rect 24814 1062 24866 1114
rect 24878 1062 24930 1114
rect 24942 1062 24994 1114
rect 1584 960 1636 1012
rect 4620 960 4672 1012
rect 7288 960 7340 1012
rect 7380 960 7432 1012
rect 15016 960 15068 1012
rect 16672 960 16724 1012
rect 16856 960 16908 1012
rect 20168 960 20220 1012
rect 2412 824 2464 876
rect 5816 824 5868 876
rect 10048 824 10100 876
rect 8484 688 8536 740
rect 9128 688 9180 740
rect 9680 688 9732 740
rect 10324 688 10376 740
rect 13636 824 13688 876
rect 23572 688 23624 740
rect 24860 688 24912 740
rect 7288 552 7340 604
rect 12532 552 12584 604
<< metal2 >>
rect 202 9840 258 10000
rect 478 9840 534 10000
rect 754 9840 810 10000
rect 1030 9840 1086 10000
rect 1306 9840 1362 10000
rect 1582 9840 1638 10000
rect 1858 9840 1914 10000
rect 2134 9840 2190 10000
rect 2410 9840 2466 10000
rect 2686 9840 2742 10000
rect 2962 9840 3018 10000
rect 3238 9840 3294 10000
rect 3514 9840 3570 10000
rect 3790 9840 3846 10000
rect 4066 9840 4122 10000
rect 4342 9840 4398 10000
rect 4618 9840 4674 10000
rect 4894 9840 4950 10000
rect 5170 9840 5226 10000
rect 5446 9840 5502 10000
rect 5722 9840 5778 10000
rect 5998 9840 6054 10000
rect 6274 9840 6330 10000
rect 6550 9840 6606 10000
rect 6826 9840 6882 10000
rect 7102 9840 7158 10000
rect 7378 9840 7434 10000
rect 7654 9840 7710 10000
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 216 6662 244 9840
rect 492 9058 520 9840
rect 492 9030 704 9058
rect 676 8566 704 9030
rect 664 8560 716 8566
rect 664 8502 716 8508
rect 204 6656 256 6662
rect 204 6598 256 6604
rect 768 6458 796 9840
rect 1044 6866 1072 9840
rect 1320 7546 1348 9840
rect 1596 8072 1624 9840
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1676 8084 1728 8090
rect 1596 8044 1676 8072
rect 1676 8026 1728 8032
rect 1780 7886 1808 9114
rect 1872 8514 1900 9840
rect 2148 9058 2176 9840
rect 2320 9240 2372 9246
rect 2320 9182 2372 9188
rect 2056 9030 2176 9058
rect 2056 8634 2084 9030
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1872 8486 2268 8514
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1950 7848 2006 7857
rect 1950 7783 2006 7792
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1964 7478 1992 7783
rect 2240 7546 2268 8486
rect 2332 7886 2360 9182
rect 2424 8090 2452 9840
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 8498 2544 9318
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2412 8084 2464 8090
rect 2700 8072 2728 9840
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2780 9308 2832 9314
rect 2780 9250 2832 9256
rect 2792 8498 2820 9250
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2780 8084 2832 8090
rect 2700 8044 2780 8072
rect 2412 8026 2464 8032
rect 2780 8026 2832 8032
rect 2884 7970 2912 9522
rect 2976 8634 3004 9840
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2700 7942 2912 7970
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2700 7478 2728 7942
rect 3160 7886 3188 8774
rect 3252 8072 3280 9840
rect 3332 8084 3384 8090
rect 3252 8044 3332 8072
rect 3332 8026 3384 8032
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 3252 7002 3280 7686
rect 3528 7206 3556 9840
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3712 9178 3740 9658
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3804 7546 3832 9840
rect 4080 8276 4108 9840
rect 4356 8634 4384 9840
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4080 8248 4292 8276
rect 3917 8188 4225 8197
rect 3917 8186 3923 8188
rect 3979 8186 4003 8188
rect 4059 8186 4083 8188
rect 4139 8186 4163 8188
rect 4219 8186 4225 8188
rect 3979 8134 3981 8186
rect 4161 8134 4163 8186
rect 3917 8132 3923 8134
rect 3979 8132 4003 8134
rect 4059 8132 4083 8134
rect 4139 8132 4163 8134
rect 4219 8132 4225 8134
rect 3917 8123 4225 8132
rect 4160 8084 4212 8090
rect 4264 8072 4292 8248
rect 4212 8044 4292 8072
rect 4160 8026 4212 8032
rect 4632 7546 4660 9840
rect 4908 8072 4936 9840
rect 5184 8634 5212 9840
rect 5460 8634 5488 9840
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5552 8498 5580 8842
rect 5736 8634 5764 9840
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 4988 8084 5040 8090
rect 4908 8044 4988 8072
rect 4988 8026 5040 8032
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5368 7546 5396 7890
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5460 7546 5488 7754
rect 5644 7546 5672 8434
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 8090 5948 8230
rect 5908 8084 5960 8090
rect 6012 8072 6040 9840
rect 6288 8090 6316 9840
rect 6092 8084 6144 8090
rect 6012 8044 6092 8072
rect 5908 8026 5960 8032
rect 6092 8026 6144 8032
rect 6276 8084 6328 8090
rect 6564 8072 6592 9840
rect 6644 9784 6696 9790
rect 6644 9726 6696 9732
rect 6656 8498 6684 9726
rect 6840 9058 6868 9840
rect 6748 9030 6868 9058
rect 6748 8634 6776 9030
rect 7116 8820 7144 9840
rect 7116 8792 7328 8820
rect 6884 8732 7192 8741
rect 6884 8730 6890 8732
rect 6946 8730 6970 8732
rect 7026 8730 7050 8732
rect 7106 8730 7130 8732
rect 7186 8730 7192 8732
rect 6946 8678 6948 8730
rect 7128 8678 7130 8730
rect 6884 8676 6890 8678
rect 6946 8676 6970 8678
rect 7026 8676 7050 8678
rect 7106 8676 7130 8678
rect 7186 8676 7192 8678
rect 6884 8667 7192 8676
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6644 8084 6696 8090
rect 6564 8044 6644 8072
rect 6276 8026 6328 8032
rect 6644 8026 6696 8032
rect 7196 8084 7248 8090
rect 7300 8072 7328 8792
rect 7392 8090 7420 9840
rect 7472 9784 7524 9790
rect 7472 9726 7524 9732
rect 7484 8498 7512 9726
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7576 8498 7604 9590
rect 7668 8634 7696 9840
rect 7852 8650 7880 9930
rect 7930 9840 7986 10000
rect 8206 9840 8262 10000
rect 8482 9840 8538 10000
rect 8758 9840 8814 10000
rect 9034 9840 9090 10000
rect 9310 9840 9366 10000
rect 9586 9840 9642 10000
rect 9862 9840 9918 10000
rect 10138 9840 10194 10000
rect 10414 9840 10470 10000
rect 10690 9840 10746 10000
rect 10966 9840 11022 10000
rect 11242 9840 11298 10000
rect 11518 9840 11574 10000
rect 11794 9840 11850 10000
rect 12070 9840 12126 10000
rect 12346 9840 12402 10000
rect 12622 9840 12678 10000
rect 12898 9840 12954 10000
rect 13174 9840 13230 10000
rect 13450 9840 13506 10000
rect 13726 9840 13782 10000
rect 14002 9840 14058 10000
rect 14278 9840 14334 10000
rect 14384 9846 14504 9874
rect 14384 9840 14412 9846
rect 7944 9432 7972 9840
rect 7944 9404 8156 9432
rect 8024 9240 8076 9246
rect 8024 9182 8076 9188
rect 7656 8628 7708 8634
rect 7852 8622 7972 8650
rect 7656 8570 7708 8576
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7248 8044 7328 8072
rect 7380 8084 7432 8090
rect 7196 8026 7248 8032
rect 7380 8026 7432 8032
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5828 7546 5856 7822
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6564 7546 6592 7754
rect 6884 7644 7192 7653
rect 6884 7642 6890 7644
rect 6946 7642 6970 7644
rect 7026 7642 7050 7644
rect 7106 7642 7130 7644
rect 7186 7642 7192 7644
rect 6946 7590 6948 7642
rect 7128 7590 7130 7642
rect 6884 7588 6890 7590
rect 6946 7588 6970 7590
rect 7026 7588 7050 7590
rect 7106 7588 7130 7590
rect 7186 7588 7192 7590
rect 6884 7579 7192 7588
rect 7378 7576 7434 7585
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 6552 7540 6604 7546
rect 7484 7546 7512 8298
rect 7378 7511 7434 7520
rect 7472 7540 7524 7546
rect 6552 7482 6604 7488
rect 5906 7440 5962 7449
rect 5906 7375 5908 7384
rect 5960 7375 5962 7384
rect 6184 7404 6236 7410
rect 5908 7346 5960 7352
rect 6184 7346 6236 7352
rect 6196 7313 6224 7346
rect 7392 7342 7420 7511
rect 7472 7482 7524 7488
rect 7576 7410 7604 8298
rect 7852 7546 7880 8502
rect 7944 7954 7972 8622
rect 8036 8566 8064 9182
rect 8128 8634 8156 9404
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8024 8560 8076 8566
rect 8220 8548 8248 9840
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8404 8838 8432 9386
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8496 8634 8524 9840
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8220 8520 8340 8548
rect 8024 8502 8076 8508
rect 8312 8090 8340 8520
rect 8392 8492 8444 8498
rect 8444 8452 8616 8480
rect 8392 8434 8444 8440
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8404 8090 8432 8230
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7380 7336 7432 7342
rect 6182 7304 6238 7313
rect 7380 7278 7432 7284
rect 6182 7239 6238 7248
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 3917 7100 4225 7109
rect 3917 7098 3923 7100
rect 3979 7098 4003 7100
rect 4059 7098 4083 7100
rect 4139 7098 4163 7100
rect 4219 7098 4225 7100
rect 3979 7046 3981 7098
rect 4161 7046 4163 7098
rect 3917 7044 3923 7046
rect 3979 7044 4003 7046
rect 4059 7044 4083 7046
rect 4139 7044 4163 7046
rect 4219 7044 4225 7046
rect 3917 7035 4225 7044
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 6288 6934 6316 7142
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 1032 6860 1084 6866
rect 1032 6802 1084 6808
rect 756 6452 808 6458
rect 756 6394 808 6400
rect 6380 6390 6408 7142
rect 7760 6730 7788 7482
rect 8128 6866 8156 7754
rect 8496 7206 8524 8230
rect 8588 7954 8616 8452
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8680 7546 8708 8842
rect 8772 8634 8800 9840
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8956 7886 8984 9454
rect 9048 8634 9076 9840
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9232 8498 9260 8774
rect 9324 8634 9352 9840
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9416 8498 9444 9046
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9600 8362 9628 9840
rect 9770 9480 9826 9489
rect 9770 9415 9826 9424
rect 9784 8430 9812 9415
rect 9876 8430 9904 9840
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9968 8566 9996 8774
rect 10152 8650 10180 9840
rect 10152 8622 10272 8650
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9864 8424 9916 8430
rect 10060 8401 10088 8434
rect 9864 8366 9916 8372
rect 10046 8392 10102 8401
rect 9588 8356 9640 8362
rect 10046 8327 10102 8336
rect 9588 8298 9640 8304
rect 9956 8288 10008 8294
rect 9692 8248 9956 8276
rect 9692 8242 9720 8248
rect 9600 8214 9720 8242
rect 9956 8230 10008 8236
rect 9600 7886 9628 8214
rect 9851 8188 10159 8197
rect 9851 8186 9857 8188
rect 9913 8186 9937 8188
rect 9993 8186 10017 8188
rect 10073 8186 10097 8188
rect 10153 8186 10159 8188
rect 9913 8134 9915 8186
rect 10095 8134 10097 8186
rect 9851 8132 9857 8134
rect 9913 8132 9937 8134
rect 9993 8132 10017 8134
rect 10073 8132 10097 8134
rect 10153 8132 10159 8134
rect 9851 8123 10159 8132
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9692 7546 9720 7958
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 7206 8708 7346
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 9784 6798 9812 7822
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10244 7698 10272 8622
rect 10428 7886 10456 9840
rect 10600 9784 10652 9790
rect 10600 9726 10652 9732
rect 10612 8498 10640 9726
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10508 7744 10560 7750
rect 10060 7585 10088 7686
rect 10244 7670 10456 7698
rect 10508 7686 10560 7692
rect 10046 7576 10102 7585
rect 10046 7511 10102 7520
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10336 7410 10364 7482
rect 10428 7410 10456 7670
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10520 7274 10548 7686
rect 10612 7274 10640 7890
rect 10704 7886 10732 9840
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10888 7750 10916 7958
rect 10980 7886 11008 9840
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8498 11192 8774
rect 11256 8514 11284 9840
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11440 8634 11468 9318
rect 11532 8922 11560 9840
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11624 9382 11652 9522
rect 11716 9489 11744 9522
rect 11702 9480 11758 9489
rect 11702 9415 11758 9424
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11808 8922 11836 9840
rect 11532 8894 11652 8922
rect 11808 8894 11928 8922
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11152 8492 11204 8498
rect 11256 8486 11468 8514
rect 11152 8434 11204 8440
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10796 7410 10824 7686
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 9851 7100 10159 7109
rect 9851 7098 9857 7100
rect 9913 7098 9937 7100
rect 9993 7098 10017 7100
rect 10073 7098 10097 7100
rect 10153 7098 10159 7100
rect 9913 7046 9915 7098
rect 10095 7046 10097 7098
rect 9851 7044 9857 7046
rect 9913 7044 9937 7046
rect 9993 7044 10017 7046
rect 10073 7044 10097 7046
rect 10153 7044 10159 7046
rect 9851 7035 10159 7044
rect 11072 7002 11100 8298
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11164 7546 11192 8026
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11348 7002 11376 8230
rect 11440 7868 11468 8486
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11532 8022 11560 8434
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11520 7880 11572 7886
rect 11440 7840 11520 7868
rect 11624 7868 11652 8894
rect 11796 7880 11848 7886
rect 11624 7840 11796 7868
rect 11520 7822 11572 7828
rect 11900 7868 11928 8894
rect 11980 8492 12032 8498
rect 12084 8480 12112 9840
rect 12360 8922 12388 9840
rect 12636 9296 12664 9840
rect 12268 8894 12388 8922
rect 12544 9268 12664 9296
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12032 8452 12112 8480
rect 11980 8434 12032 8440
rect 12176 7954 12204 8570
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12072 7880 12124 7886
rect 11900 7840 12072 7868
rect 11796 7822 11848 7828
rect 12268 7868 12296 8894
rect 12544 8498 12572 9268
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12636 8634 12664 9114
rect 12912 8922 12940 9840
rect 13188 9058 13216 9840
rect 13188 9030 13308 9058
rect 12912 8894 13216 8922
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12728 8498 12756 8774
rect 12818 8732 13126 8741
rect 12818 8730 12824 8732
rect 12880 8730 12904 8732
rect 12960 8730 12984 8732
rect 13040 8730 13064 8732
rect 13120 8730 13126 8732
rect 12880 8678 12882 8730
rect 13062 8678 13064 8730
rect 12818 8676 12824 8678
rect 12880 8676 12904 8678
rect 12960 8676 12984 8678
rect 13040 8676 13064 8678
rect 13120 8676 13126 8678
rect 12818 8667 13126 8676
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12440 8424 12492 8430
rect 12808 8424 12860 8430
rect 12492 8372 12808 8378
rect 12440 8366 12860 8372
rect 12990 8392 13046 8401
rect 12452 8350 12848 8366
rect 12990 8327 13046 8336
rect 13004 8090 13032 8327
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13188 7886 13216 8894
rect 12348 7880 12400 7886
rect 12268 7840 12348 7868
rect 12072 7822 12124 7828
rect 12348 7822 12400 7828
rect 13176 7880 13228 7886
rect 13280 7868 13308 9030
rect 13360 8492 13412 8498
rect 13464 8480 13492 9840
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13556 8498 13584 9386
rect 13412 8452 13492 8480
rect 13544 8492 13596 8498
rect 13360 8434 13412 8440
rect 13544 8434 13596 8440
rect 13636 8492 13688 8498
rect 13740 8480 13768 9840
rect 13912 9308 13964 9314
rect 13912 9250 13964 9256
rect 13924 8634 13952 9250
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14016 8566 14044 9840
rect 14292 9812 14412 9840
rect 14096 9784 14148 9790
rect 14096 9726 14148 9732
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13688 8452 13768 8480
rect 13636 8434 13688 8440
rect 14108 8090 14136 9726
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 8634 14228 9318
rect 14476 8634 14504 9846
rect 14554 9840 14610 10000
rect 14830 9840 14886 10000
rect 15016 9852 15068 9858
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14200 8090 14228 8434
rect 14476 8362 14504 8434
rect 14568 8430 14596 9840
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14384 8242 14412 8298
rect 14752 8294 14780 8774
rect 14556 8288 14608 8294
rect 14384 8236 14556 8242
rect 14384 8230 14608 8236
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14384 8214 14596 8230
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14844 7886 14872 9840
rect 15106 9840 15162 10000
rect 15382 9840 15438 10000
rect 15658 9840 15714 10000
rect 15934 9840 15990 10000
rect 16210 9840 16266 10000
rect 16486 9840 16542 10000
rect 16762 9840 16818 10000
rect 17038 9840 17094 10000
rect 17314 9840 17370 10000
rect 17590 9840 17646 10000
rect 17866 9840 17922 10000
rect 18142 9840 18198 10000
rect 18418 9840 18474 10000
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 15016 9794 15068 9800
rect 15028 8294 15056 9794
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 13452 7880 13504 7886
rect 13280 7840 13452 7868
rect 13176 7822 13228 7828
rect 13452 7822 13504 7828
rect 14832 7880 14884 7886
rect 15120 7868 15148 9840
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15212 8634 15240 9658
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15212 8090 15240 8434
rect 15396 8362 15424 9840
rect 15672 8922 15700 9840
rect 15580 8894 15700 8922
rect 15948 8922 15976 9840
rect 15844 8900 15896 8906
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15384 7880 15436 7886
rect 15120 7840 15384 7868
rect 14832 7822 14884 7828
rect 15488 7857 15516 8570
rect 15384 7822 15436 7828
rect 15474 7848 15530 7857
rect 15474 7783 15530 7792
rect 15580 7800 15608 8894
rect 15948 8894 16160 8922
rect 15844 8842 15896 8848
rect 15856 8634 15884 8842
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15672 8090 15700 8434
rect 15785 8188 16093 8197
rect 15785 8186 15791 8188
rect 15847 8186 15871 8188
rect 15927 8186 15951 8188
rect 16007 8186 16031 8188
rect 16087 8186 16093 8188
rect 15847 8134 15849 8186
rect 16029 8134 16031 8186
rect 15785 8132 15791 8134
rect 15847 8132 15871 8134
rect 15927 8132 15951 8134
rect 16007 8132 16031 8134
rect 16087 8132 16093 8134
rect 15785 8123 16093 8132
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 16132 7886 16160 8894
rect 16224 7954 16252 9840
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16316 8634 16344 9454
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 15660 7812 15712 7818
rect 15580 7772 15660 7800
rect 15660 7754 15712 7760
rect 12818 7644 13126 7653
rect 12818 7642 12824 7644
rect 12880 7642 12904 7644
rect 12960 7642 12984 7644
rect 13040 7642 13064 7644
rect 13120 7642 13126 7644
rect 12880 7590 12882 7642
rect 13062 7590 13064 7642
rect 12818 7588 12824 7590
rect 12880 7588 12904 7590
rect 12960 7588 12984 7590
rect 13040 7588 13064 7590
rect 13120 7588 13126 7590
rect 12818 7579 13126 7588
rect 15785 7100 16093 7109
rect 15785 7098 15791 7100
rect 15847 7098 15871 7100
rect 15927 7098 15951 7100
rect 16007 7098 16031 7100
rect 16087 7098 16093 7100
rect 15847 7046 15849 7098
rect 16029 7046 16031 7098
rect 15785 7044 15791 7046
rect 15847 7044 15871 7046
rect 15927 7044 15951 7046
rect 16007 7044 16031 7046
rect 16087 7044 16093 7046
rect 15785 7035 16093 7044
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 6884 6556 7192 6565
rect 6884 6554 6890 6556
rect 6946 6554 6970 6556
rect 7026 6554 7050 6556
rect 7106 6554 7130 6556
rect 7186 6554 7192 6556
rect 6946 6502 6948 6554
rect 7128 6502 7130 6554
rect 6884 6500 6890 6502
rect 6946 6500 6970 6502
rect 7026 6500 7050 6502
rect 7106 6500 7130 6502
rect 7186 6500 7192 6502
rect 6884 6491 7192 6500
rect 12818 6556 13126 6565
rect 12818 6554 12824 6556
rect 12880 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13126 6556
rect 12880 6502 12882 6554
rect 13062 6502 13064 6554
rect 12818 6500 12824 6502
rect 12880 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13126 6502
rect 12818 6491 13126 6500
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 9851 6012 10159 6021
rect 9851 6010 9857 6012
rect 9913 6010 9937 6012
rect 9993 6010 10017 6012
rect 10073 6010 10097 6012
rect 10153 6010 10159 6012
rect 9913 5958 9915 6010
rect 10095 5958 10097 6010
rect 9851 5956 9857 5958
rect 9913 5956 9937 5958
rect 9993 5956 10017 5958
rect 10073 5956 10097 5958
rect 10153 5956 10159 5958
rect 9851 5947 10159 5956
rect 15785 6012 16093 6021
rect 15785 6010 15791 6012
rect 15847 6010 15871 6012
rect 15927 6010 15951 6012
rect 16007 6010 16031 6012
rect 16087 6010 16093 6012
rect 15847 5958 15849 6010
rect 16029 5958 16031 6010
rect 15785 5956 15791 5958
rect 15847 5956 15871 5958
rect 15927 5956 15951 5958
rect 16007 5956 16031 5958
rect 16087 5956 16093 5958
rect 15785 5947 16093 5956
rect 6884 5468 7192 5477
rect 6884 5466 6890 5468
rect 6946 5466 6970 5468
rect 7026 5466 7050 5468
rect 7106 5466 7130 5468
rect 7186 5466 7192 5468
rect 6946 5414 6948 5466
rect 7128 5414 7130 5466
rect 6884 5412 6890 5414
rect 6946 5412 6970 5414
rect 7026 5412 7050 5414
rect 7106 5412 7130 5414
rect 7186 5412 7192 5414
rect 6884 5403 7192 5412
rect 12818 5468 13126 5477
rect 12818 5466 12824 5468
rect 12880 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13126 5468
rect 12880 5414 12882 5466
rect 13062 5414 13064 5466
rect 12818 5412 12824 5414
rect 12880 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13126 5414
rect 12818 5403 13126 5412
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 9851 4924 10159 4933
rect 9851 4922 9857 4924
rect 9913 4922 9937 4924
rect 9993 4922 10017 4924
rect 10073 4922 10097 4924
rect 10153 4922 10159 4924
rect 9913 4870 9915 4922
rect 10095 4870 10097 4922
rect 9851 4868 9857 4870
rect 9913 4868 9937 4870
rect 9993 4868 10017 4870
rect 10073 4868 10097 4870
rect 10153 4868 10159 4870
rect 9851 4859 10159 4868
rect 15785 4924 16093 4933
rect 15785 4922 15791 4924
rect 15847 4922 15871 4924
rect 15927 4922 15951 4924
rect 16007 4922 16031 4924
rect 16087 4922 16093 4924
rect 15847 4870 15849 4922
rect 16029 4870 16031 4922
rect 15785 4868 15791 4870
rect 15847 4868 15871 4870
rect 15927 4868 15951 4870
rect 16007 4868 16031 4870
rect 16087 4868 16093 4870
rect 15785 4859 16093 4868
rect 6884 4380 7192 4389
rect 6884 4378 6890 4380
rect 6946 4378 6970 4380
rect 7026 4378 7050 4380
rect 7106 4378 7130 4380
rect 7186 4378 7192 4380
rect 6946 4326 6948 4378
rect 7128 4326 7130 4378
rect 6884 4324 6890 4326
rect 6946 4324 6970 4326
rect 7026 4324 7050 4326
rect 7106 4324 7130 4326
rect 7186 4324 7192 4326
rect 6884 4315 7192 4324
rect 12818 4380 13126 4389
rect 12818 4378 12824 4380
rect 12880 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13126 4380
rect 12880 4326 12882 4378
rect 13062 4326 13064 4378
rect 12818 4324 12824 4326
rect 12880 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13126 4326
rect 12818 4315 13126 4324
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 9851 3836 10159 3845
rect 9851 3834 9857 3836
rect 9913 3834 9937 3836
rect 9993 3834 10017 3836
rect 10073 3834 10097 3836
rect 10153 3834 10159 3836
rect 9913 3782 9915 3834
rect 10095 3782 10097 3834
rect 9851 3780 9857 3782
rect 9913 3780 9937 3782
rect 9993 3780 10017 3782
rect 10073 3780 10097 3782
rect 10153 3780 10159 3782
rect 9851 3771 10159 3780
rect 15785 3836 16093 3845
rect 15785 3834 15791 3836
rect 15847 3834 15871 3836
rect 15927 3834 15951 3836
rect 16007 3834 16031 3836
rect 16087 3834 16093 3836
rect 15847 3782 15849 3834
rect 16029 3782 16031 3834
rect 15785 3780 15791 3782
rect 15847 3780 15871 3782
rect 15927 3780 15951 3782
rect 16007 3780 16031 3782
rect 16087 3780 16093 3782
rect 15785 3771 16093 3780
rect 6884 3292 7192 3301
rect 6884 3290 6890 3292
rect 6946 3290 6970 3292
rect 7026 3290 7050 3292
rect 7106 3290 7130 3292
rect 7186 3290 7192 3292
rect 6946 3238 6948 3290
rect 7128 3238 7130 3290
rect 6884 3236 6890 3238
rect 6946 3236 6970 3238
rect 7026 3236 7050 3238
rect 7106 3236 7130 3238
rect 7186 3236 7192 3238
rect 6884 3227 7192 3236
rect 12818 3292 13126 3301
rect 12818 3290 12824 3292
rect 12880 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13126 3292
rect 12880 3238 12882 3290
rect 13062 3238 13064 3290
rect 12818 3236 12824 3238
rect 12880 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13126 3238
rect 12818 3227 13126 3236
rect 16408 2774 16436 8570
rect 16500 8022 16528 9840
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16684 8634 16712 9046
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16684 7750 16712 8366
rect 16776 7818 16804 9840
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16960 8634 16988 8978
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16868 8090 16896 8434
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 17052 7954 17080 9840
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17236 8634 17264 8910
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17236 8022 17264 8366
rect 17328 8022 17356 9840
rect 17500 9240 17552 9246
rect 17500 9182 17552 9188
rect 17512 8634 17540 9182
rect 17604 8634 17632 9840
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17880 8537 17908 9840
rect 17866 8528 17922 8537
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17776 8492 17828 8498
rect 17866 8463 17922 8472
rect 17776 8434 17828 8440
rect 17420 8090 17448 8434
rect 17788 8090 17816 8434
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 8090 17908 8230
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 18156 7886 18184 9840
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18248 8362 18276 9590
rect 18432 8378 18460 9840
rect 18524 8514 18552 9862
rect 18616 8634 18644 9930
rect 18694 9840 18750 10000
rect 18970 9840 19026 10000
rect 19246 9840 19302 10000
rect 19522 9840 19578 10000
rect 19798 9840 19854 10000
rect 20074 9840 20130 10000
rect 20350 9840 20406 10000
rect 20626 9840 20682 10000
rect 20902 9840 20958 10000
rect 21178 9840 21234 10000
rect 21454 9840 21510 10000
rect 21730 9840 21786 10000
rect 22006 9840 22062 10000
rect 22282 9840 22338 10000
rect 22558 9840 22614 10000
rect 22834 9840 22890 10000
rect 23110 9840 23166 10000
rect 23386 9840 23442 10000
rect 23662 9840 23718 10000
rect 23938 9840 23994 10000
rect 24214 9840 24270 10000
rect 24490 9840 24546 10000
rect 24766 9840 24822 10000
rect 25042 9840 25098 10000
rect 25318 9840 25374 10000
rect 25594 9840 25650 10000
rect 18708 9178 18736 9840
rect 18984 9194 19012 9840
rect 18696 9172 18748 9178
rect 18984 9166 19196 9194
rect 18696 9114 18748 9120
rect 18752 8732 19060 8741
rect 18752 8730 18758 8732
rect 18814 8730 18838 8732
rect 18894 8730 18918 8732
rect 18974 8730 18998 8732
rect 19054 8730 19060 8732
rect 18814 8678 18816 8730
rect 18996 8678 18998 8730
rect 18752 8676 18758 8678
rect 18814 8676 18838 8678
rect 18894 8676 18918 8678
rect 18974 8676 18998 8678
rect 19054 8676 19060 8678
rect 18752 8667 19060 8676
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 19168 8566 19196 9166
rect 18972 8560 19024 8566
rect 18970 8528 18972 8537
rect 19156 8560 19208 8566
rect 19024 8528 19026 8537
rect 18524 8486 18828 8514
rect 18604 8424 18656 8430
rect 18432 8372 18604 8378
rect 18432 8366 18656 8372
rect 18236 8356 18288 8362
rect 18432 8350 18644 8366
rect 18236 8298 18288 8304
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 8090 18644 8230
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18800 8022 18828 8486
rect 18880 8492 18932 8498
rect 19156 8502 19208 8508
rect 18970 8463 19026 8472
rect 18880 8434 18932 8440
rect 18892 8090 18920 8434
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 19168 7886 19196 8230
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 19156 7880 19208 7886
rect 19260 7868 19288 9840
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 8090 19380 8230
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19340 7880 19392 7886
rect 19260 7840 19340 7868
rect 19156 7822 19208 7828
rect 19536 7868 19564 9840
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19720 8498 19748 9114
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19616 7880 19668 7886
rect 19536 7840 19616 7868
rect 19340 7822 19392 7828
rect 19812 7868 19840 9840
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19996 8634 20024 9522
rect 20088 8634 20116 9840
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20076 8628 20128 8634
rect 20364 8616 20392 9840
rect 20536 8628 20588 8634
rect 20364 8588 20536 8616
rect 20076 8570 20128 8576
rect 20640 8616 20668 9840
rect 20916 8786 20944 9840
rect 20916 8758 21036 8786
rect 20904 8628 20956 8634
rect 20640 8588 20904 8616
rect 20536 8570 20588 8576
rect 20904 8570 20956 8576
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 19892 7880 19944 7886
rect 19812 7840 19892 7868
rect 19616 7822 19668 7828
rect 19892 7822 19944 7828
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17512 5914 17540 6258
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 9851 2748 10159 2757
rect 9851 2746 9857 2748
rect 9913 2746 9937 2748
rect 9993 2746 10017 2748
rect 10073 2746 10097 2748
rect 10153 2746 10159 2748
rect 9913 2694 9915 2746
rect 10095 2694 10097 2746
rect 9851 2692 9857 2694
rect 9913 2692 9937 2694
rect 9993 2692 10017 2694
rect 10073 2692 10097 2694
rect 10153 2692 10159 2694
rect 9851 2683 10159 2692
rect 15785 2748 16093 2757
rect 15785 2746 15791 2748
rect 15847 2746 15871 2748
rect 15927 2746 15951 2748
rect 16007 2746 16031 2748
rect 16087 2746 16093 2748
rect 15847 2694 15849 2746
rect 16029 2694 16031 2746
rect 15785 2692 15791 2694
rect 15847 2692 15871 2694
rect 15927 2692 15951 2694
rect 16007 2692 16031 2694
rect 16087 2692 16093 2694
rect 15785 2683 16093 2692
rect 16316 2746 16436 2774
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 11702 2544 11758 2553
rect 11702 2479 11758 2488
rect 10230 2408 10286 2417
rect 10230 2343 10286 2352
rect 6884 2204 7192 2213
rect 6884 2202 6890 2204
rect 6946 2202 6970 2204
rect 7026 2202 7050 2204
rect 7106 2202 7130 2204
rect 7186 2202 7192 2204
rect 6946 2150 6948 2202
rect 7128 2150 7130 2202
rect 6884 2148 6890 2150
rect 6946 2148 6970 2150
rect 7026 2148 7050 2150
rect 7106 2148 7130 2150
rect 7186 2148 7192 2150
rect 6884 2139 7192 2148
rect 10244 2106 10272 2343
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10612 2106 10640 2246
rect 11716 2106 11744 2479
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 12818 2204 13126 2213
rect 12818 2202 12824 2204
rect 12880 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13126 2204
rect 12880 2150 12882 2202
rect 13062 2150 13064 2202
rect 12818 2148 12824 2150
rect 12880 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13126 2150
rect 12818 2139 13126 2148
rect 13740 2106 13768 2382
rect 13832 2106 13860 2586
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15120 2106 15148 2518
rect 9128 2100 9180 2106
rect 9128 2042 9180 2048
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10600 2100 10652 2106
rect 10600 2042 10652 2048
rect 11704 2100 11756 2106
rect 11704 2042 11756 2048
rect 13728 2100 13780 2106
rect 13728 2042 13780 2048
rect 13820 2100 13872 2106
rect 13820 2042 13872 2048
rect 15108 2100 15160 2106
rect 15108 2042 15160 2048
rect 9140 2009 9168 2042
rect 9126 2000 9182 2009
rect 7748 1964 7800 1970
rect 7748 1906 7800 1912
rect 8944 1964 8996 1970
rect 16316 1970 16344 2746
rect 9126 1935 9182 1944
rect 9772 1964 9824 1970
rect 8944 1906 8996 1912
rect 9772 1906 9824 1912
rect 10416 1964 10468 1970
rect 10416 1906 10468 1912
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 12624 1964 12676 1970
rect 12624 1906 12676 1912
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 13912 1964 13964 1970
rect 13912 1906 13964 1912
rect 14924 1964 14976 1970
rect 14924 1906 14976 1912
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 3917 1660 4225 1669
rect 3917 1658 3923 1660
rect 3979 1658 4003 1660
rect 4059 1658 4083 1660
rect 4139 1658 4163 1660
rect 4219 1658 4225 1660
rect 3979 1606 3981 1658
rect 4161 1606 4163 1658
rect 3917 1604 3923 1606
rect 3979 1604 4003 1606
rect 4059 1604 4083 1606
rect 4139 1604 4163 1606
rect 4219 1604 4225 1606
rect 3917 1595 4225 1604
rect 7760 1562 7788 1906
rect 7930 1864 7986 1873
rect 7930 1799 7932 1808
rect 7984 1799 7986 1808
rect 7932 1770 7984 1776
rect 8956 1562 8984 1906
rect 9784 1562 9812 1906
rect 9851 1660 10159 1669
rect 9851 1658 9857 1660
rect 9913 1658 9937 1660
rect 9993 1658 10017 1660
rect 10073 1658 10097 1660
rect 10153 1658 10159 1660
rect 9913 1606 9915 1658
rect 10095 1606 10097 1658
rect 9851 1604 9857 1606
rect 9913 1604 9937 1606
rect 9993 1604 10017 1606
rect 10073 1604 10097 1606
rect 10153 1604 10159 1606
rect 9851 1595 10159 1604
rect 10428 1562 10456 1906
rect 11532 1562 11560 1906
rect 7748 1556 7800 1562
rect 7748 1498 7800 1504
rect 8944 1556 8996 1562
rect 8944 1498 8996 1504
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 10416 1556 10468 1562
rect 10416 1498 10468 1504
rect 11520 1556 11572 1562
rect 11520 1498 11572 1504
rect 940 1352 992 1358
rect 940 1294 992 1300
rect 2228 1352 2280 1358
rect 2228 1294 2280 1300
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 6000 1352 6052 1358
rect 7656 1352 7708 1358
rect 6000 1294 6052 1300
rect 7484 1312 7656 1340
rect 952 160 980 1294
rect 1584 1216 1636 1222
rect 1584 1158 1636 1164
rect 1596 1018 1624 1158
rect 1584 1012 1636 1018
rect 1584 954 1636 960
rect 938 0 994 160
rect 2134 82 2190 160
rect 2240 82 2268 1294
rect 2412 1216 2464 1222
rect 2412 1158 2464 1164
rect 2424 882 2452 1158
rect 2412 876 2464 882
rect 2412 818 2464 824
rect 2134 54 2268 82
rect 3330 82 3386 160
rect 3436 82 3464 1294
rect 4620 1216 4672 1222
rect 4620 1158 4672 1164
rect 4632 1018 4660 1158
rect 4620 1012 4672 1018
rect 4620 954 4672 960
rect 3330 54 3464 82
rect 4526 82 4582 160
rect 4816 82 4844 1294
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 5828 882 5856 1158
rect 5816 876 5868 882
rect 5816 818 5868 824
rect 4526 54 4844 82
rect 5722 82 5778 160
rect 6012 82 6040 1294
rect 7380 1216 7432 1222
rect 7380 1158 7432 1164
rect 6884 1116 7192 1125
rect 6884 1114 6890 1116
rect 6946 1114 6970 1116
rect 7026 1114 7050 1116
rect 7106 1114 7130 1116
rect 7186 1114 7192 1116
rect 6946 1062 6948 1114
rect 7128 1062 7130 1114
rect 6884 1060 6890 1062
rect 6946 1060 6970 1062
rect 7026 1060 7050 1062
rect 7106 1060 7130 1062
rect 7186 1060 7192 1062
rect 6884 1051 7192 1060
rect 7392 1018 7420 1158
rect 7288 1012 7340 1018
rect 7288 954 7340 960
rect 7380 1012 7432 1018
rect 7380 954 7432 960
rect 7300 610 7328 954
rect 7288 604 7340 610
rect 7288 546 7340 552
rect 5722 54 6040 82
rect 6918 82 6974 160
rect 7484 82 7512 1312
rect 7656 1294 7708 1300
rect 9128 1352 9180 1358
rect 9128 1294 9180 1300
rect 10048 1352 10100 1358
rect 10048 1294 10100 1300
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 10784 1352 10836 1358
rect 10784 1294 10836 1300
rect 11980 1352 12032 1358
rect 11980 1294 12032 1300
rect 12532 1352 12584 1358
rect 12532 1294 12584 1300
rect 9140 746 9168 1294
rect 10060 882 10088 1294
rect 10048 876 10100 882
rect 10048 818 10100 824
rect 10336 746 10364 1294
rect 8484 740 8536 746
rect 8484 682 8536 688
rect 9128 740 9180 746
rect 9128 682 9180 688
rect 9680 740 9732 746
rect 9680 682 9732 688
rect 10324 740 10376 746
rect 10324 682 10376 688
rect 6918 54 7512 82
rect 8114 82 8170 160
rect 8496 82 8524 682
rect 8114 54 8524 82
rect 9310 82 9366 160
rect 9692 82 9720 682
rect 9310 54 9720 82
rect 10506 82 10562 160
rect 10796 82 10824 1294
rect 10506 54 10824 82
rect 11702 82 11758 160
rect 11992 82 12020 1294
rect 12544 610 12572 1294
rect 12636 1222 12664 1906
rect 12912 1562 12940 1906
rect 13648 1562 13676 1906
rect 13924 1562 13952 1906
rect 14936 1562 14964 1906
rect 12900 1556 12952 1562
rect 12900 1498 12952 1504
rect 13636 1556 13688 1562
rect 13636 1498 13688 1504
rect 13912 1556 13964 1562
rect 13912 1498 13964 1504
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 13268 1420 13320 1426
rect 13268 1362 13320 1368
rect 12624 1216 12676 1222
rect 12624 1158 12676 1164
rect 12818 1116 13126 1125
rect 12818 1114 12824 1116
rect 12880 1114 12904 1116
rect 12960 1114 12984 1116
rect 13040 1114 13064 1116
rect 13120 1114 13126 1116
rect 12880 1062 12882 1114
rect 13062 1062 13064 1114
rect 12818 1060 12824 1062
rect 12880 1060 12904 1062
rect 12960 1060 12984 1062
rect 13040 1060 13064 1062
rect 13120 1060 13126 1062
rect 12818 1051 13126 1060
rect 12532 604 12584 610
rect 12532 546 12584 552
rect 12912 190 13032 218
rect 12912 160 12940 190
rect 11702 54 12020 82
rect 2134 0 2190 54
rect 3330 0 3386 54
rect 4526 0 4582 54
rect 5722 0 5778 54
rect 6918 0 6974 54
rect 8114 0 8170 54
rect 9310 0 9366 54
rect 10506 0 10562 54
rect 11702 0 11758 54
rect 12898 0 12954 160
rect 13004 82 13032 190
rect 13280 82 13308 1362
rect 15396 1358 15424 1906
rect 15785 1660 16093 1669
rect 15785 1658 15791 1660
rect 15847 1658 15871 1660
rect 15927 1658 15951 1660
rect 16007 1658 16031 1660
rect 16087 1658 16093 1660
rect 15847 1606 15849 1658
rect 16029 1606 16031 1658
rect 15785 1604 15791 1606
rect 15847 1604 15871 1606
rect 15927 1604 15951 1606
rect 16007 1604 16031 1606
rect 16087 1604 16093 1606
rect 15785 1595 16093 1604
rect 16132 1562 16160 1906
rect 16120 1556 16172 1562
rect 16120 1498 16172 1504
rect 16960 1358 16988 5646
rect 17788 2106 17816 7482
rect 18064 7002 18092 7686
rect 18752 7644 19060 7653
rect 18752 7642 18758 7644
rect 18814 7642 18838 7644
rect 18894 7642 18918 7644
rect 18974 7642 18998 7644
rect 19054 7642 19060 7644
rect 18814 7590 18816 7642
rect 18996 7590 18998 7642
rect 18752 7588 18758 7590
rect 18814 7588 18838 7590
rect 18894 7588 18918 7590
rect 18974 7588 18998 7590
rect 19054 7588 19060 7590
rect 18752 7579 19060 7588
rect 19536 7313 19564 7686
rect 19812 7478 19840 7686
rect 19800 7472 19852 7478
rect 20088 7449 20116 7686
rect 19800 7414 19852 7420
rect 20074 7440 20130 7449
rect 20074 7375 20130 7384
rect 19522 7304 19578 7313
rect 19522 7239 19578 7248
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18752 6556 19060 6565
rect 18752 6554 18758 6556
rect 18814 6554 18838 6556
rect 18894 6554 18918 6556
rect 18974 6554 18998 6556
rect 19054 6554 19060 6556
rect 18814 6502 18816 6554
rect 18996 6502 18998 6554
rect 18752 6500 18758 6502
rect 18814 6500 18838 6502
rect 18894 6500 18918 6502
rect 18974 6500 18998 6502
rect 19054 6500 19060 6502
rect 18752 6491 19060 6500
rect 18752 5468 19060 5477
rect 18752 5466 18758 5468
rect 18814 5466 18838 5468
rect 18894 5466 18918 5468
rect 18974 5466 18998 5468
rect 19054 5466 19060 5468
rect 18814 5414 18816 5466
rect 18996 5414 18998 5466
rect 18752 5412 18758 5414
rect 18814 5412 18838 5414
rect 18894 5412 18918 5414
rect 18974 5412 18998 5414
rect 19054 5412 19060 5414
rect 18752 5403 19060 5412
rect 18752 4380 19060 4389
rect 18752 4378 18758 4380
rect 18814 4378 18838 4380
rect 18894 4378 18918 4380
rect 18974 4378 18998 4380
rect 19054 4378 19060 4380
rect 18814 4326 18816 4378
rect 18996 4326 18998 4378
rect 18752 4324 18758 4326
rect 18814 4324 18838 4326
rect 18894 4324 18918 4326
rect 18974 4324 18998 4326
rect 19054 4324 19060 4326
rect 18752 4315 19060 4324
rect 18752 3292 19060 3301
rect 18752 3290 18758 3292
rect 18814 3290 18838 3292
rect 18894 3290 18918 3292
rect 18974 3290 18998 3292
rect 19054 3290 19060 3292
rect 18814 3238 18816 3290
rect 18996 3238 18998 3290
rect 18752 3236 18758 3238
rect 18814 3236 18838 3238
rect 18894 3236 18918 3238
rect 18974 3236 18998 3238
rect 19054 3236 19060 3238
rect 18752 3227 19060 3236
rect 18752 2204 19060 2213
rect 18752 2202 18758 2204
rect 18814 2202 18838 2204
rect 18894 2202 18918 2204
rect 18974 2202 18998 2204
rect 19054 2202 19060 2204
rect 18814 2150 18816 2202
rect 18996 2150 18998 2202
rect 18752 2148 18758 2150
rect 18814 2148 18838 2150
rect 18894 2148 18918 2150
rect 18974 2148 18998 2150
rect 19054 2148 19060 2150
rect 18752 2139 19060 2148
rect 17776 2100 17828 2106
rect 17776 2042 17828 2048
rect 18604 1964 18656 1970
rect 18604 1906 18656 1912
rect 18616 1562 18644 1906
rect 18604 1556 18656 1562
rect 18604 1498 18656 1504
rect 13636 1352 13688 1358
rect 13636 1294 13688 1300
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 15016 1352 15068 1358
rect 15016 1294 15068 1300
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15568 1352 15620 1358
rect 15568 1294 15620 1300
rect 16672 1352 16724 1358
rect 16672 1294 16724 1300
rect 16948 1352 17000 1358
rect 17132 1352 17184 1358
rect 16948 1294 17000 1300
rect 17052 1312 17132 1340
rect 13648 882 13676 1294
rect 13636 876 13688 882
rect 13636 818 13688 824
rect 13004 54 13308 82
rect 14094 82 14150 160
rect 14384 82 14412 1294
rect 15028 1018 15056 1294
rect 15016 1012 15068 1018
rect 15016 954 15068 960
rect 14094 54 14412 82
rect 15290 82 15346 160
rect 15580 82 15608 1294
rect 16684 1018 16712 1294
rect 16856 1216 16908 1222
rect 16856 1158 16908 1164
rect 16868 1018 16896 1158
rect 16672 1012 16724 1018
rect 16672 954 16724 960
rect 16856 1012 16908 1018
rect 16856 954 16908 960
rect 15290 54 15608 82
rect 16486 82 16542 160
rect 17052 82 17080 1312
rect 17132 1294 17184 1300
rect 17960 1352 18012 1358
rect 19432 1352 19484 1358
rect 17960 1294 18012 1300
rect 19352 1312 19432 1340
rect 16486 54 17080 82
rect 17682 82 17738 160
rect 17972 82 18000 1294
rect 18752 1116 19060 1125
rect 18752 1114 18758 1116
rect 18814 1114 18838 1116
rect 18894 1114 18918 1116
rect 18974 1114 18998 1116
rect 19054 1114 19060 1116
rect 18814 1062 18816 1114
rect 18996 1062 18998 1114
rect 18752 1060 18758 1062
rect 18814 1060 18838 1062
rect 18894 1060 18918 1062
rect 18974 1060 18998 1062
rect 19054 1060 19060 1062
rect 18752 1051 19060 1060
rect 17682 54 18000 82
rect 18878 82 18934 160
rect 19352 82 19380 1312
rect 19432 1294 19484 1300
rect 20180 1018 20208 8434
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20732 1970 20760 7346
rect 20536 1964 20588 1970
rect 20536 1906 20588 1912
rect 20720 1964 20772 1970
rect 20720 1906 20772 1912
rect 20548 1562 20576 1906
rect 20824 1766 20852 8434
rect 21008 8430 21036 8758
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21192 8090 21220 9840
rect 21468 8616 21496 9840
rect 21744 9110 21772 9840
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21548 8628 21600 8634
rect 21468 8588 21548 8616
rect 21548 8570 21600 8576
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20916 2310 20944 7822
rect 21284 2446 21312 8434
rect 22020 8276 22048 9840
rect 22296 8786 22324 9840
rect 22572 8888 22600 9840
rect 22572 8860 22692 8888
rect 22296 8758 22600 8786
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22020 8248 22140 8276
rect 21719 8188 22027 8197
rect 21719 8186 21725 8188
rect 21781 8186 21805 8188
rect 21861 8186 21885 8188
rect 21941 8186 21965 8188
rect 22021 8186 22027 8188
rect 21781 8134 21783 8186
rect 21963 8134 21965 8186
rect 21719 8132 21725 8134
rect 21781 8132 21805 8134
rect 21861 8132 21885 8134
rect 21941 8132 21965 8134
rect 22021 8132 22027 8134
rect 21719 8123 22027 8132
rect 21916 7812 21968 7818
rect 21916 7754 21968 7760
rect 21928 7546 21956 7754
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21719 7100 22027 7109
rect 21719 7098 21725 7100
rect 21781 7098 21805 7100
rect 21861 7098 21885 7100
rect 21941 7098 21965 7100
rect 22021 7098 22027 7100
rect 21781 7046 21783 7098
rect 21963 7046 21965 7098
rect 21719 7044 21725 7046
rect 21781 7044 21805 7046
rect 21861 7044 21885 7046
rect 21941 7044 21965 7046
rect 22021 7044 22027 7046
rect 21719 7035 22027 7044
rect 22112 7002 22140 8248
rect 22296 7698 22324 8434
rect 22480 7970 22508 8434
rect 22572 8090 22600 8758
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22664 7970 22692 8860
rect 22848 8090 22876 9840
rect 22928 9104 22980 9110
rect 22928 9046 22980 9052
rect 22940 8634 22968 9046
rect 23124 8634 23152 9840
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22204 7670 22324 7698
rect 22388 7942 22508 7970
rect 22572 7942 22692 7970
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21719 6012 22027 6021
rect 21719 6010 21725 6012
rect 21781 6010 21805 6012
rect 21861 6010 21885 6012
rect 21941 6010 21965 6012
rect 22021 6010 22027 6012
rect 21781 5958 21783 6010
rect 21963 5958 21965 6010
rect 21719 5956 21725 5958
rect 21781 5956 21805 5958
rect 21861 5956 21885 5958
rect 21941 5956 21965 5958
rect 22021 5956 22027 5958
rect 21719 5947 22027 5956
rect 21719 4924 22027 4933
rect 21719 4922 21725 4924
rect 21781 4922 21805 4924
rect 21861 4922 21885 4924
rect 21941 4922 21965 4924
rect 22021 4922 22027 4924
rect 21781 4870 21783 4922
rect 21963 4870 21965 4922
rect 21719 4868 21725 4870
rect 21781 4868 21805 4870
rect 21861 4868 21885 4870
rect 21941 4868 21965 4870
rect 22021 4868 22027 4870
rect 21719 4859 22027 4868
rect 21719 3836 22027 3845
rect 21719 3834 21725 3836
rect 21781 3834 21805 3836
rect 21861 3834 21885 3836
rect 21941 3834 21965 3836
rect 22021 3834 22027 3836
rect 21781 3782 21783 3834
rect 21963 3782 21965 3834
rect 21719 3780 21725 3782
rect 21781 3780 21805 3782
rect 21861 3780 21885 3782
rect 21941 3780 21965 3782
rect 22021 3780 22027 3782
rect 21719 3771 22027 3780
rect 21719 2748 22027 2757
rect 21719 2746 21725 2748
rect 21781 2746 21805 2748
rect 21861 2746 21885 2748
rect 21941 2746 21965 2748
rect 22021 2746 22027 2748
rect 21781 2694 21783 2746
rect 21963 2694 21965 2746
rect 21719 2692 21725 2694
rect 21781 2692 21805 2694
rect 21861 2692 21885 2694
rect 21941 2692 21965 2694
rect 22021 2692 22027 2694
rect 21719 2683 22027 2692
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 22112 2106 22140 6734
rect 22100 2100 22152 2106
rect 22100 2042 22152 2048
rect 22204 1873 22232 7670
rect 22388 6914 22416 7942
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22296 6886 22416 6914
rect 22296 2281 22324 6886
rect 22480 2553 22508 7754
rect 22572 7546 22600 7942
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22664 2650 22692 7754
rect 22940 2650 22968 8434
rect 23400 8090 23428 9840
rect 23676 8090 23704 9840
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23848 7812 23900 7818
rect 23848 7754 23900 7760
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23020 6724 23072 6730
rect 23020 6666 23072 6672
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 22466 2544 22522 2553
rect 22466 2479 22522 2488
rect 22376 2440 22428 2446
rect 23032 2417 23060 6666
rect 22376 2382 22428 2388
rect 23018 2408 23074 2417
rect 22282 2272 22338 2281
rect 22282 2207 22338 2216
rect 22388 2106 22416 2382
rect 23018 2343 23074 2352
rect 23124 2106 23152 7346
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 23308 2378 23336 7278
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23296 2372 23348 2378
rect 23296 2314 23348 2320
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 23112 2100 23164 2106
rect 23112 2042 23164 2048
rect 22284 1964 22336 1970
rect 22284 1906 22336 1912
rect 22560 1964 22612 1970
rect 22560 1906 22612 1912
rect 22190 1864 22246 1873
rect 22190 1799 22246 1808
rect 20812 1760 20864 1766
rect 20812 1702 20864 1708
rect 21719 1660 22027 1669
rect 21719 1658 21725 1660
rect 21781 1658 21805 1660
rect 21861 1658 21885 1660
rect 21941 1658 21965 1660
rect 22021 1658 22027 1660
rect 21781 1606 21783 1658
rect 21963 1606 21965 1658
rect 21719 1604 21725 1606
rect 21781 1604 21805 1606
rect 21861 1604 21885 1606
rect 21941 1604 21965 1606
rect 22021 1604 22027 1606
rect 21719 1595 22027 1604
rect 22296 1562 22324 1906
rect 22572 1562 22600 1906
rect 23400 1834 23428 6326
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23492 1834 23520 6258
rect 23676 2446 23704 7346
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23768 2106 23796 7686
rect 23860 6118 23888 7754
rect 23952 6458 23980 9840
rect 24228 7546 24256 9840
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24504 6458 24532 9840
rect 24780 8888 24808 9840
rect 24596 8860 24808 8888
rect 24596 6866 24624 8860
rect 24686 8732 24994 8741
rect 24686 8730 24692 8732
rect 24748 8730 24772 8732
rect 24828 8730 24852 8732
rect 24908 8730 24932 8732
rect 24988 8730 24994 8732
rect 24748 8678 24750 8730
rect 24930 8678 24932 8730
rect 24686 8676 24692 8678
rect 24748 8676 24772 8678
rect 24828 8676 24852 8678
rect 24908 8676 24932 8678
rect 24988 8676 24994 8678
rect 24686 8667 24994 8676
rect 24686 7644 24994 7653
rect 24686 7642 24692 7644
rect 24748 7642 24772 7644
rect 24828 7642 24852 7644
rect 24908 7642 24932 7644
rect 24988 7642 24994 7644
rect 24748 7590 24750 7642
rect 24930 7590 24932 7642
rect 24686 7588 24692 7590
rect 24748 7588 24772 7590
rect 24828 7588 24852 7590
rect 24908 7588 24932 7590
rect 24988 7588 24994 7590
rect 24686 7579 24994 7588
rect 25056 7342 25084 9840
rect 25332 7546 25360 9840
rect 25608 7886 25636 9840
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24686 6556 24994 6565
rect 24686 6554 24692 6556
rect 24748 6554 24772 6556
rect 24828 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 24994 6556
rect 24748 6502 24750 6554
rect 24930 6502 24932 6554
rect 24686 6500 24692 6502
rect 24748 6500 24772 6502
rect 24828 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 24994 6502
rect 24686 6491 24994 6500
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 24686 5468 24994 5477
rect 24686 5466 24692 5468
rect 24748 5466 24772 5468
rect 24828 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 24994 5468
rect 24748 5414 24750 5466
rect 24930 5414 24932 5466
rect 24686 5412 24692 5414
rect 24748 5412 24772 5414
rect 24828 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 24994 5414
rect 24686 5403 24994 5412
rect 24686 4380 24994 4389
rect 24686 4378 24692 4380
rect 24748 4378 24772 4380
rect 24828 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 24994 4380
rect 24748 4326 24750 4378
rect 24930 4326 24932 4378
rect 24686 4324 24692 4326
rect 24748 4324 24772 4326
rect 24828 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 24994 4326
rect 24686 4315 24994 4324
rect 24686 3292 24994 3301
rect 24686 3290 24692 3292
rect 24748 3290 24772 3292
rect 24828 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 24994 3292
rect 24748 3238 24750 3290
rect 24930 3238 24932 3290
rect 24686 3236 24692 3238
rect 24748 3236 24772 3238
rect 24828 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 24994 3238
rect 24686 3227 24994 3236
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 24136 2106 24164 2314
rect 24686 2204 24994 2213
rect 24686 2202 24692 2204
rect 24748 2202 24772 2204
rect 24828 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 24994 2204
rect 24748 2150 24750 2202
rect 24930 2150 24932 2202
rect 24686 2148 24692 2150
rect 24748 2148 24772 2150
rect 24828 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 24994 2150
rect 24686 2139 24994 2148
rect 23756 2100 23808 2106
rect 23756 2042 23808 2048
rect 24124 2100 24176 2106
rect 24124 2042 24176 2048
rect 23572 1964 23624 1970
rect 23572 1906 23624 1912
rect 24032 1964 24084 1970
rect 24032 1906 24084 1912
rect 24308 1964 24360 1970
rect 24308 1906 24360 1912
rect 23388 1828 23440 1834
rect 23388 1770 23440 1776
rect 23480 1828 23532 1834
rect 23480 1770 23532 1776
rect 23584 1562 23612 1906
rect 20536 1556 20588 1562
rect 20536 1498 20588 1504
rect 22284 1556 22336 1562
rect 22284 1498 22336 1504
rect 22560 1556 22612 1562
rect 22560 1498 22612 1504
rect 23572 1556 23624 1562
rect 23572 1498 23624 1504
rect 24044 1494 24072 1906
rect 24320 1562 24348 1906
rect 24308 1556 24360 1562
rect 24308 1498 24360 1504
rect 24032 1488 24084 1494
rect 24032 1430 24084 1436
rect 20352 1352 20404 1358
rect 20352 1294 20404 1300
rect 21548 1352 21600 1358
rect 21548 1294 21600 1300
rect 22744 1352 22796 1358
rect 22744 1294 22796 1300
rect 23572 1352 23624 1358
rect 23572 1294 23624 1300
rect 24216 1352 24268 1358
rect 24216 1294 24268 1300
rect 20168 1012 20220 1018
rect 20168 954 20220 960
rect 18878 54 19380 82
rect 20074 82 20130 160
rect 20364 82 20392 1294
rect 20074 54 20392 82
rect 21270 82 21326 160
rect 21560 82 21588 1294
rect 21270 54 21588 82
rect 22466 82 22522 160
rect 22756 82 22784 1294
rect 23584 746 23612 1294
rect 23572 740 23624 746
rect 23572 682 23624 688
rect 24228 218 24256 1294
rect 24686 1116 24994 1125
rect 24686 1114 24692 1116
rect 24748 1114 24772 1116
rect 24828 1114 24852 1116
rect 24908 1114 24932 1116
rect 24988 1114 24994 1116
rect 24748 1062 24750 1114
rect 24930 1062 24932 1114
rect 24686 1060 24692 1062
rect 24748 1060 24772 1062
rect 24828 1060 24852 1062
rect 24908 1060 24932 1062
rect 24988 1060 24994 1062
rect 24686 1051 24994 1060
rect 24860 740 24912 746
rect 24860 682 24912 688
rect 23676 190 23796 218
rect 23676 160 23704 190
rect 22466 54 22784 82
rect 14094 0 14150 54
rect 15290 0 15346 54
rect 16486 0 16542 54
rect 17682 0 17738 54
rect 18878 0 18934 54
rect 20074 0 20130 54
rect 21270 0 21326 54
rect 22466 0 22522 54
rect 23662 0 23718 160
rect 23768 82 23796 190
rect 24136 190 24256 218
rect 24136 82 24164 190
rect 24872 160 24900 682
rect 23768 54 24164 82
rect 24858 0 24914 160
<< via2 >>
rect 1950 7792 2006 7848
rect 3923 8186 3979 8188
rect 4003 8186 4059 8188
rect 4083 8186 4139 8188
rect 4163 8186 4219 8188
rect 3923 8134 3969 8186
rect 3969 8134 3979 8186
rect 4003 8134 4033 8186
rect 4033 8134 4045 8186
rect 4045 8134 4059 8186
rect 4083 8134 4097 8186
rect 4097 8134 4109 8186
rect 4109 8134 4139 8186
rect 4163 8134 4173 8186
rect 4173 8134 4219 8186
rect 3923 8132 3979 8134
rect 4003 8132 4059 8134
rect 4083 8132 4139 8134
rect 4163 8132 4219 8134
rect 6890 8730 6946 8732
rect 6970 8730 7026 8732
rect 7050 8730 7106 8732
rect 7130 8730 7186 8732
rect 6890 8678 6936 8730
rect 6936 8678 6946 8730
rect 6970 8678 7000 8730
rect 7000 8678 7012 8730
rect 7012 8678 7026 8730
rect 7050 8678 7064 8730
rect 7064 8678 7076 8730
rect 7076 8678 7106 8730
rect 7130 8678 7140 8730
rect 7140 8678 7186 8730
rect 6890 8676 6946 8678
rect 6970 8676 7026 8678
rect 7050 8676 7106 8678
rect 7130 8676 7186 8678
rect 6890 7642 6946 7644
rect 6970 7642 7026 7644
rect 7050 7642 7106 7644
rect 7130 7642 7186 7644
rect 6890 7590 6936 7642
rect 6936 7590 6946 7642
rect 6970 7590 7000 7642
rect 7000 7590 7012 7642
rect 7012 7590 7026 7642
rect 7050 7590 7064 7642
rect 7064 7590 7076 7642
rect 7076 7590 7106 7642
rect 7130 7590 7140 7642
rect 7140 7590 7186 7642
rect 6890 7588 6946 7590
rect 6970 7588 7026 7590
rect 7050 7588 7106 7590
rect 7130 7588 7186 7590
rect 7378 7520 7434 7576
rect 5906 7404 5962 7440
rect 5906 7384 5908 7404
rect 5908 7384 5960 7404
rect 5960 7384 5962 7404
rect 6182 7248 6238 7304
rect 3923 7098 3979 7100
rect 4003 7098 4059 7100
rect 4083 7098 4139 7100
rect 4163 7098 4219 7100
rect 3923 7046 3969 7098
rect 3969 7046 3979 7098
rect 4003 7046 4033 7098
rect 4033 7046 4045 7098
rect 4045 7046 4059 7098
rect 4083 7046 4097 7098
rect 4097 7046 4109 7098
rect 4109 7046 4139 7098
rect 4163 7046 4173 7098
rect 4173 7046 4219 7098
rect 3923 7044 3979 7046
rect 4003 7044 4059 7046
rect 4083 7044 4139 7046
rect 4163 7044 4219 7046
rect 9770 9424 9826 9480
rect 10046 8336 10102 8392
rect 9857 8186 9913 8188
rect 9937 8186 9993 8188
rect 10017 8186 10073 8188
rect 10097 8186 10153 8188
rect 9857 8134 9903 8186
rect 9903 8134 9913 8186
rect 9937 8134 9967 8186
rect 9967 8134 9979 8186
rect 9979 8134 9993 8186
rect 10017 8134 10031 8186
rect 10031 8134 10043 8186
rect 10043 8134 10073 8186
rect 10097 8134 10107 8186
rect 10107 8134 10153 8186
rect 9857 8132 9913 8134
rect 9937 8132 9993 8134
rect 10017 8132 10073 8134
rect 10097 8132 10153 8134
rect 10046 7520 10102 7576
rect 11702 9424 11758 9480
rect 9857 7098 9913 7100
rect 9937 7098 9993 7100
rect 10017 7098 10073 7100
rect 10097 7098 10153 7100
rect 9857 7046 9903 7098
rect 9903 7046 9913 7098
rect 9937 7046 9967 7098
rect 9967 7046 9979 7098
rect 9979 7046 9993 7098
rect 10017 7046 10031 7098
rect 10031 7046 10043 7098
rect 10043 7046 10073 7098
rect 10097 7046 10107 7098
rect 10107 7046 10153 7098
rect 9857 7044 9913 7046
rect 9937 7044 9993 7046
rect 10017 7044 10073 7046
rect 10097 7044 10153 7046
rect 12824 8730 12880 8732
rect 12904 8730 12960 8732
rect 12984 8730 13040 8732
rect 13064 8730 13120 8732
rect 12824 8678 12870 8730
rect 12870 8678 12880 8730
rect 12904 8678 12934 8730
rect 12934 8678 12946 8730
rect 12946 8678 12960 8730
rect 12984 8678 12998 8730
rect 12998 8678 13010 8730
rect 13010 8678 13040 8730
rect 13064 8678 13074 8730
rect 13074 8678 13120 8730
rect 12824 8676 12880 8678
rect 12904 8676 12960 8678
rect 12984 8676 13040 8678
rect 13064 8676 13120 8678
rect 12990 8336 13046 8392
rect 15474 7792 15530 7848
rect 15791 8186 15847 8188
rect 15871 8186 15927 8188
rect 15951 8186 16007 8188
rect 16031 8186 16087 8188
rect 15791 8134 15837 8186
rect 15837 8134 15847 8186
rect 15871 8134 15901 8186
rect 15901 8134 15913 8186
rect 15913 8134 15927 8186
rect 15951 8134 15965 8186
rect 15965 8134 15977 8186
rect 15977 8134 16007 8186
rect 16031 8134 16041 8186
rect 16041 8134 16087 8186
rect 15791 8132 15847 8134
rect 15871 8132 15927 8134
rect 15951 8132 16007 8134
rect 16031 8132 16087 8134
rect 12824 7642 12880 7644
rect 12904 7642 12960 7644
rect 12984 7642 13040 7644
rect 13064 7642 13120 7644
rect 12824 7590 12870 7642
rect 12870 7590 12880 7642
rect 12904 7590 12934 7642
rect 12934 7590 12946 7642
rect 12946 7590 12960 7642
rect 12984 7590 12998 7642
rect 12998 7590 13010 7642
rect 13010 7590 13040 7642
rect 13064 7590 13074 7642
rect 13074 7590 13120 7642
rect 12824 7588 12880 7590
rect 12904 7588 12960 7590
rect 12984 7588 13040 7590
rect 13064 7588 13120 7590
rect 15791 7098 15847 7100
rect 15871 7098 15927 7100
rect 15951 7098 16007 7100
rect 16031 7098 16087 7100
rect 15791 7046 15837 7098
rect 15837 7046 15847 7098
rect 15871 7046 15901 7098
rect 15901 7046 15913 7098
rect 15913 7046 15927 7098
rect 15951 7046 15965 7098
rect 15965 7046 15977 7098
rect 15977 7046 16007 7098
rect 16031 7046 16041 7098
rect 16041 7046 16087 7098
rect 15791 7044 15847 7046
rect 15871 7044 15927 7046
rect 15951 7044 16007 7046
rect 16031 7044 16087 7046
rect 6890 6554 6946 6556
rect 6970 6554 7026 6556
rect 7050 6554 7106 6556
rect 7130 6554 7186 6556
rect 6890 6502 6936 6554
rect 6936 6502 6946 6554
rect 6970 6502 7000 6554
rect 7000 6502 7012 6554
rect 7012 6502 7026 6554
rect 7050 6502 7064 6554
rect 7064 6502 7076 6554
rect 7076 6502 7106 6554
rect 7130 6502 7140 6554
rect 7140 6502 7186 6554
rect 6890 6500 6946 6502
rect 6970 6500 7026 6502
rect 7050 6500 7106 6502
rect 7130 6500 7186 6502
rect 12824 6554 12880 6556
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 12824 6502 12870 6554
rect 12870 6502 12880 6554
rect 12904 6502 12934 6554
rect 12934 6502 12946 6554
rect 12946 6502 12960 6554
rect 12984 6502 12998 6554
rect 12998 6502 13010 6554
rect 13010 6502 13040 6554
rect 13064 6502 13074 6554
rect 13074 6502 13120 6554
rect 12824 6500 12880 6502
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 9857 6010 9913 6012
rect 9937 6010 9993 6012
rect 10017 6010 10073 6012
rect 10097 6010 10153 6012
rect 9857 5958 9903 6010
rect 9903 5958 9913 6010
rect 9937 5958 9967 6010
rect 9967 5958 9979 6010
rect 9979 5958 9993 6010
rect 10017 5958 10031 6010
rect 10031 5958 10043 6010
rect 10043 5958 10073 6010
rect 10097 5958 10107 6010
rect 10107 5958 10153 6010
rect 9857 5956 9913 5958
rect 9937 5956 9993 5958
rect 10017 5956 10073 5958
rect 10097 5956 10153 5958
rect 15791 6010 15847 6012
rect 15871 6010 15927 6012
rect 15951 6010 16007 6012
rect 16031 6010 16087 6012
rect 15791 5958 15837 6010
rect 15837 5958 15847 6010
rect 15871 5958 15901 6010
rect 15901 5958 15913 6010
rect 15913 5958 15927 6010
rect 15951 5958 15965 6010
rect 15965 5958 15977 6010
rect 15977 5958 16007 6010
rect 16031 5958 16041 6010
rect 16041 5958 16087 6010
rect 15791 5956 15847 5958
rect 15871 5956 15927 5958
rect 15951 5956 16007 5958
rect 16031 5956 16087 5958
rect 6890 5466 6946 5468
rect 6970 5466 7026 5468
rect 7050 5466 7106 5468
rect 7130 5466 7186 5468
rect 6890 5414 6936 5466
rect 6936 5414 6946 5466
rect 6970 5414 7000 5466
rect 7000 5414 7012 5466
rect 7012 5414 7026 5466
rect 7050 5414 7064 5466
rect 7064 5414 7076 5466
rect 7076 5414 7106 5466
rect 7130 5414 7140 5466
rect 7140 5414 7186 5466
rect 6890 5412 6946 5414
rect 6970 5412 7026 5414
rect 7050 5412 7106 5414
rect 7130 5412 7186 5414
rect 12824 5466 12880 5468
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 12824 5414 12870 5466
rect 12870 5414 12880 5466
rect 12904 5414 12934 5466
rect 12934 5414 12946 5466
rect 12946 5414 12960 5466
rect 12984 5414 12998 5466
rect 12998 5414 13010 5466
rect 13010 5414 13040 5466
rect 13064 5414 13074 5466
rect 13074 5414 13120 5466
rect 12824 5412 12880 5414
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 9857 4922 9913 4924
rect 9937 4922 9993 4924
rect 10017 4922 10073 4924
rect 10097 4922 10153 4924
rect 9857 4870 9903 4922
rect 9903 4870 9913 4922
rect 9937 4870 9967 4922
rect 9967 4870 9979 4922
rect 9979 4870 9993 4922
rect 10017 4870 10031 4922
rect 10031 4870 10043 4922
rect 10043 4870 10073 4922
rect 10097 4870 10107 4922
rect 10107 4870 10153 4922
rect 9857 4868 9913 4870
rect 9937 4868 9993 4870
rect 10017 4868 10073 4870
rect 10097 4868 10153 4870
rect 15791 4922 15847 4924
rect 15871 4922 15927 4924
rect 15951 4922 16007 4924
rect 16031 4922 16087 4924
rect 15791 4870 15837 4922
rect 15837 4870 15847 4922
rect 15871 4870 15901 4922
rect 15901 4870 15913 4922
rect 15913 4870 15927 4922
rect 15951 4870 15965 4922
rect 15965 4870 15977 4922
rect 15977 4870 16007 4922
rect 16031 4870 16041 4922
rect 16041 4870 16087 4922
rect 15791 4868 15847 4870
rect 15871 4868 15927 4870
rect 15951 4868 16007 4870
rect 16031 4868 16087 4870
rect 6890 4378 6946 4380
rect 6970 4378 7026 4380
rect 7050 4378 7106 4380
rect 7130 4378 7186 4380
rect 6890 4326 6936 4378
rect 6936 4326 6946 4378
rect 6970 4326 7000 4378
rect 7000 4326 7012 4378
rect 7012 4326 7026 4378
rect 7050 4326 7064 4378
rect 7064 4326 7076 4378
rect 7076 4326 7106 4378
rect 7130 4326 7140 4378
rect 7140 4326 7186 4378
rect 6890 4324 6946 4326
rect 6970 4324 7026 4326
rect 7050 4324 7106 4326
rect 7130 4324 7186 4326
rect 12824 4378 12880 4380
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 12824 4326 12870 4378
rect 12870 4326 12880 4378
rect 12904 4326 12934 4378
rect 12934 4326 12946 4378
rect 12946 4326 12960 4378
rect 12984 4326 12998 4378
rect 12998 4326 13010 4378
rect 13010 4326 13040 4378
rect 13064 4326 13074 4378
rect 13074 4326 13120 4378
rect 12824 4324 12880 4326
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 9857 3834 9913 3836
rect 9937 3834 9993 3836
rect 10017 3834 10073 3836
rect 10097 3834 10153 3836
rect 9857 3782 9903 3834
rect 9903 3782 9913 3834
rect 9937 3782 9967 3834
rect 9967 3782 9979 3834
rect 9979 3782 9993 3834
rect 10017 3782 10031 3834
rect 10031 3782 10043 3834
rect 10043 3782 10073 3834
rect 10097 3782 10107 3834
rect 10107 3782 10153 3834
rect 9857 3780 9913 3782
rect 9937 3780 9993 3782
rect 10017 3780 10073 3782
rect 10097 3780 10153 3782
rect 15791 3834 15847 3836
rect 15871 3834 15927 3836
rect 15951 3834 16007 3836
rect 16031 3834 16087 3836
rect 15791 3782 15837 3834
rect 15837 3782 15847 3834
rect 15871 3782 15901 3834
rect 15901 3782 15913 3834
rect 15913 3782 15927 3834
rect 15951 3782 15965 3834
rect 15965 3782 15977 3834
rect 15977 3782 16007 3834
rect 16031 3782 16041 3834
rect 16041 3782 16087 3834
rect 15791 3780 15847 3782
rect 15871 3780 15927 3782
rect 15951 3780 16007 3782
rect 16031 3780 16087 3782
rect 6890 3290 6946 3292
rect 6970 3290 7026 3292
rect 7050 3290 7106 3292
rect 7130 3290 7186 3292
rect 6890 3238 6936 3290
rect 6936 3238 6946 3290
rect 6970 3238 7000 3290
rect 7000 3238 7012 3290
rect 7012 3238 7026 3290
rect 7050 3238 7064 3290
rect 7064 3238 7076 3290
rect 7076 3238 7106 3290
rect 7130 3238 7140 3290
rect 7140 3238 7186 3290
rect 6890 3236 6946 3238
rect 6970 3236 7026 3238
rect 7050 3236 7106 3238
rect 7130 3236 7186 3238
rect 12824 3290 12880 3292
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 12824 3238 12870 3290
rect 12870 3238 12880 3290
rect 12904 3238 12934 3290
rect 12934 3238 12946 3290
rect 12946 3238 12960 3290
rect 12984 3238 12998 3290
rect 12998 3238 13010 3290
rect 13010 3238 13040 3290
rect 13064 3238 13074 3290
rect 13074 3238 13120 3290
rect 12824 3236 12880 3238
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 17866 8472 17922 8528
rect 18758 8730 18814 8732
rect 18838 8730 18894 8732
rect 18918 8730 18974 8732
rect 18998 8730 19054 8732
rect 18758 8678 18804 8730
rect 18804 8678 18814 8730
rect 18838 8678 18868 8730
rect 18868 8678 18880 8730
rect 18880 8678 18894 8730
rect 18918 8678 18932 8730
rect 18932 8678 18944 8730
rect 18944 8678 18974 8730
rect 18998 8678 19008 8730
rect 19008 8678 19054 8730
rect 18758 8676 18814 8678
rect 18838 8676 18894 8678
rect 18918 8676 18974 8678
rect 18998 8676 19054 8678
rect 18970 8508 18972 8528
rect 18972 8508 19024 8528
rect 19024 8508 19026 8528
rect 18970 8472 19026 8508
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 9857 2746 9913 2748
rect 9937 2746 9993 2748
rect 10017 2746 10073 2748
rect 10097 2746 10153 2748
rect 9857 2694 9903 2746
rect 9903 2694 9913 2746
rect 9937 2694 9967 2746
rect 9967 2694 9979 2746
rect 9979 2694 9993 2746
rect 10017 2694 10031 2746
rect 10031 2694 10043 2746
rect 10043 2694 10073 2746
rect 10097 2694 10107 2746
rect 10107 2694 10153 2746
rect 9857 2692 9913 2694
rect 9937 2692 9993 2694
rect 10017 2692 10073 2694
rect 10097 2692 10153 2694
rect 15791 2746 15847 2748
rect 15871 2746 15927 2748
rect 15951 2746 16007 2748
rect 16031 2746 16087 2748
rect 15791 2694 15837 2746
rect 15837 2694 15847 2746
rect 15871 2694 15901 2746
rect 15901 2694 15913 2746
rect 15913 2694 15927 2746
rect 15951 2694 15965 2746
rect 15965 2694 15977 2746
rect 15977 2694 16007 2746
rect 16031 2694 16041 2746
rect 16041 2694 16087 2746
rect 15791 2692 15847 2694
rect 15871 2692 15927 2694
rect 15951 2692 16007 2694
rect 16031 2692 16087 2694
rect 11702 2488 11758 2544
rect 10230 2352 10286 2408
rect 6890 2202 6946 2204
rect 6970 2202 7026 2204
rect 7050 2202 7106 2204
rect 7130 2202 7186 2204
rect 6890 2150 6936 2202
rect 6936 2150 6946 2202
rect 6970 2150 7000 2202
rect 7000 2150 7012 2202
rect 7012 2150 7026 2202
rect 7050 2150 7064 2202
rect 7064 2150 7076 2202
rect 7076 2150 7106 2202
rect 7130 2150 7140 2202
rect 7140 2150 7186 2202
rect 6890 2148 6946 2150
rect 6970 2148 7026 2150
rect 7050 2148 7106 2150
rect 7130 2148 7186 2150
rect 12824 2202 12880 2204
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 12824 2150 12870 2202
rect 12870 2150 12880 2202
rect 12904 2150 12934 2202
rect 12934 2150 12946 2202
rect 12946 2150 12960 2202
rect 12984 2150 12998 2202
rect 12998 2150 13010 2202
rect 13010 2150 13040 2202
rect 13064 2150 13074 2202
rect 13074 2150 13120 2202
rect 12824 2148 12880 2150
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 9126 1944 9182 2000
rect 3923 1658 3979 1660
rect 4003 1658 4059 1660
rect 4083 1658 4139 1660
rect 4163 1658 4219 1660
rect 3923 1606 3969 1658
rect 3969 1606 3979 1658
rect 4003 1606 4033 1658
rect 4033 1606 4045 1658
rect 4045 1606 4059 1658
rect 4083 1606 4097 1658
rect 4097 1606 4109 1658
rect 4109 1606 4139 1658
rect 4163 1606 4173 1658
rect 4173 1606 4219 1658
rect 3923 1604 3979 1606
rect 4003 1604 4059 1606
rect 4083 1604 4139 1606
rect 4163 1604 4219 1606
rect 7930 1828 7986 1864
rect 7930 1808 7932 1828
rect 7932 1808 7984 1828
rect 7984 1808 7986 1828
rect 9857 1658 9913 1660
rect 9937 1658 9993 1660
rect 10017 1658 10073 1660
rect 10097 1658 10153 1660
rect 9857 1606 9903 1658
rect 9903 1606 9913 1658
rect 9937 1606 9967 1658
rect 9967 1606 9979 1658
rect 9979 1606 9993 1658
rect 10017 1606 10031 1658
rect 10031 1606 10043 1658
rect 10043 1606 10073 1658
rect 10097 1606 10107 1658
rect 10107 1606 10153 1658
rect 9857 1604 9913 1606
rect 9937 1604 9993 1606
rect 10017 1604 10073 1606
rect 10097 1604 10153 1606
rect 6890 1114 6946 1116
rect 6970 1114 7026 1116
rect 7050 1114 7106 1116
rect 7130 1114 7186 1116
rect 6890 1062 6936 1114
rect 6936 1062 6946 1114
rect 6970 1062 7000 1114
rect 7000 1062 7012 1114
rect 7012 1062 7026 1114
rect 7050 1062 7064 1114
rect 7064 1062 7076 1114
rect 7076 1062 7106 1114
rect 7130 1062 7140 1114
rect 7140 1062 7186 1114
rect 6890 1060 6946 1062
rect 6970 1060 7026 1062
rect 7050 1060 7106 1062
rect 7130 1060 7186 1062
rect 12824 1114 12880 1116
rect 12904 1114 12960 1116
rect 12984 1114 13040 1116
rect 13064 1114 13120 1116
rect 12824 1062 12870 1114
rect 12870 1062 12880 1114
rect 12904 1062 12934 1114
rect 12934 1062 12946 1114
rect 12946 1062 12960 1114
rect 12984 1062 12998 1114
rect 12998 1062 13010 1114
rect 13010 1062 13040 1114
rect 13064 1062 13074 1114
rect 13074 1062 13120 1114
rect 12824 1060 12880 1062
rect 12904 1060 12960 1062
rect 12984 1060 13040 1062
rect 13064 1060 13120 1062
rect 15791 1658 15847 1660
rect 15871 1658 15927 1660
rect 15951 1658 16007 1660
rect 16031 1658 16087 1660
rect 15791 1606 15837 1658
rect 15837 1606 15847 1658
rect 15871 1606 15901 1658
rect 15901 1606 15913 1658
rect 15913 1606 15927 1658
rect 15951 1606 15965 1658
rect 15965 1606 15977 1658
rect 15977 1606 16007 1658
rect 16031 1606 16041 1658
rect 16041 1606 16087 1658
rect 15791 1604 15847 1606
rect 15871 1604 15927 1606
rect 15951 1604 16007 1606
rect 16031 1604 16087 1606
rect 18758 7642 18814 7644
rect 18838 7642 18894 7644
rect 18918 7642 18974 7644
rect 18998 7642 19054 7644
rect 18758 7590 18804 7642
rect 18804 7590 18814 7642
rect 18838 7590 18868 7642
rect 18868 7590 18880 7642
rect 18880 7590 18894 7642
rect 18918 7590 18932 7642
rect 18932 7590 18944 7642
rect 18944 7590 18974 7642
rect 18998 7590 19008 7642
rect 19008 7590 19054 7642
rect 18758 7588 18814 7590
rect 18838 7588 18894 7590
rect 18918 7588 18974 7590
rect 18998 7588 19054 7590
rect 20074 7384 20130 7440
rect 19522 7248 19578 7304
rect 18758 6554 18814 6556
rect 18838 6554 18894 6556
rect 18918 6554 18974 6556
rect 18998 6554 19054 6556
rect 18758 6502 18804 6554
rect 18804 6502 18814 6554
rect 18838 6502 18868 6554
rect 18868 6502 18880 6554
rect 18880 6502 18894 6554
rect 18918 6502 18932 6554
rect 18932 6502 18944 6554
rect 18944 6502 18974 6554
rect 18998 6502 19008 6554
rect 19008 6502 19054 6554
rect 18758 6500 18814 6502
rect 18838 6500 18894 6502
rect 18918 6500 18974 6502
rect 18998 6500 19054 6502
rect 18758 5466 18814 5468
rect 18838 5466 18894 5468
rect 18918 5466 18974 5468
rect 18998 5466 19054 5468
rect 18758 5414 18804 5466
rect 18804 5414 18814 5466
rect 18838 5414 18868 5466
rect 18868 5414 18880 5466
rect 18880 5414 18894 5466
rect 18918 5414 18932 5466
rect 18932 5414 18944 5466
rect 18944 5414 18974 5466
rect 18998 5414 19008 5466
rect 19008 5414 19054 5466
rect 18758 5412 18814 5414
rect 18838 5412 18894 5414
rect 18918 5412 18974 5414
rect 18998 5412 19054 5414
rect 18758 4378 18814 4380
rect 18838 4378 18894 4380
rect 18918 4378 18974 4380
rect 18998 4378 19054 4380
rect 18758 4326 18804 4378
rect 18804 4326 18814 4378
rect 18838 4326 18868 4378
rect 18868 4326 18880 4378
rect 18880 4326 18894 4378
rect 18918 4326 18932 4378
rect 18932 4326 18944 4378
rect 18944 4326 18974 4378
rect 18998 4326 19008 4378
rect 19008 4326 19054 4378
rect 18758 4324 18814 4326
rect 18838 4324 18894 4326
rect 18918 4324 18974 4326
rect 18998 4324 19054 4326
rect 18758 3290 18814 3292
rect 18838 3290 18894 3292
rect 18918 3290 18974 3292
rect 18998 3290 19054 3292
rect 18758 3238 18804 3290
rect 18804 3238 18814 3290
rect 18838 3238 18868 3290
rect 18868 3238 18880 3290
rect 18880 3238 18894 3290
rect 18918 3238 18932 3290
rect 18932 3238 18944 3290
rect 18944 3238 18974 3290
rect 18998 3238 19008 3290
rect 19008 3238 19054 3290
rect 18758 3236 18814 3238
rect 18838 3236 18894 3238
rect 18918 3236 18974 3238
rect 18998 3236 19054 3238
rect 18758 2202 18814 2204
rect 18838 2202 18894 2204
rect 18918 2202 18974 2204
rect 18998 2202 19054 2204
rect 18758 2150 18804 2202
rect 18804 2150 18814 2202
rect 18838 2150 18868 2202
rect 18868 2150 18880 2202
rect 18880 2150 18894 2202
rect 18918 2150 18932 2202
rect 18932 2150 18944 2202
rect 18944 2150 18974 2202
rect 18998 2150 19008 2202
rect 19008 2150 19054 2202
rect 18758 2148 18814 2150
rect 18838 2148 18894 2150
rect 18918 2148 18974 2150
rect 18998 2148 19054 2150
rect 18758 1114 18814 1116
rect 18838 1114 18894 1116
rect 18918 1114 18974 1116
rect 18998 1114 19054 1116
rect 18758 1062 18804 1114
rect 18804 1062 18814 1114
rect 18838 1062 18868 1114
rect 18868 1062 18880 1114
rect 18880 1062 18894 1114
rect 18918 1062 18932 1114
rect 18932 1062 18944 1114
rect 18944 1062 18974 1114
rect 18998 1062 19008 1114
rect 19008 1062 19054 1114
rect 18758 1060 18814 1062
rect 18838 1060 18894 1062
rect 18918 1060 18974 1062
rect 18998 1060 19054 1062
rect 21725 8186 21781 8188
rect 21805 8186 21861 8188
rect 21885 8186 21941 8188
rect 21965 8186 22021 8188
rect 21725 8134 21771 8186
rect 21771 8134 21781 8186
rect 21805 8134 21835 8186
rect 21835 8134 21847 8186
rect 21847 8134 21861 8186
rect 21885 8134 21899 8186
rect 21899 8134 21911 8186
rect 21911 8134 21941 8186
rect 21965 8134 21975 8186
rect 21975 8134 22021 8186
rect 21725 8132 21781 8134
rect 21805 8132 21861 8134
rect 21885 8132 21941 8134
rect 21965 8132 22021 8134
rect 21725 7098 21781 7100
rect 21805 7098 21861 7100
rect 21885 7098 21941 7100
rect 21965 7098 22021 7100
rect 21725 7046 21771 7098
rect 21771 7046 21781 7098
rect 21805 7046 21835 7098
rect 21835 7046 21847 7098
rect 21847 7046 21861 7098
rect 21885 7046 21899 7098
rect 21899 7046 21911 7098
rect 21911 7046 21941 7098
rect 21965 7046 21975 7098
rect 21975 7046 22021 7098
rect 21725 7044 21781 7046
rect 21805 7044 21861 7046
rect 21885 7044 21941 7046
rect 21965 7044 22021 7046
rect 21725 6010 21781 6012
rect 21805 6010 21861 6012
rect 21885 6010 21941 6012
rect 21965 6010 22021 6012
rect 21725 5958 21771 6010
rect 21771 5958 21781 6010
rect 21805 5958 21835 6010
rect 21835 5958 21847 6010
rect 21847 5958 21861 6010
rect 21885 5958 21899 6010
rect 21899 5958 21911 6010
rect 21911 5958 21941 6010
rect 21965 5958 21975 6010
rect 21975 5958 22021 6010
rect 21725 5956 21781 5958
rect 21805 5956 21861 5958
rect 21885 5956 21941 5958
rect 21965 5956 22021 5958
rect 21725 4922 21781 4924
rect 21805 4922 21861 4924
rect 21885 4922 21941 4924
rect 21965 4922 22021 4924
rect 21725 4870 21771 4922
rect 21771 4870 21781 4922
rect 21805 4870 21835 4922
rect 21835 4870 21847 4922
rect 21847 4870 21861 4922
rect 21885 4870 21899 4922
rect 21899 4870 21911 4922
rect 21911 4870 21941 4922
rect 21965 4870 21975 4922
rect 21975 4870 22021 4922
rect 21725 4868 21781 4870
rect 21805 4868 21861 4870
rect 21885 4868 21941 4870
rect 21965 4868 22021 4870
rect 21725 3834 21781 3836
rect 21805 3834 21861 3836
rect 21885 3834 21941 3836
rect 21965 3834 22021 3836
rect 21725 3782 21771 3834
rect 21771 3782 21781 3834
rect 21805 3782 21835 3834
rect 21835 3782 21847 3834
rect 21847 3782 21861 3834
rect 21885 3782 21899 3834
rect 21899 3782 21911 3834
rect 21911 3782 21941 3834
rect 21965 3782 21975 3834
rect 21975 3782 22021 3834
rect 21725 3780 21781 3782
rect 21805 3780 21861 3782
rect 21885 3780 21941 3782
rect 21965 3780 22021 3782
rect 21725 2746 21781 2748
rect 21805 2746 21861 2748
rect 21885 2746 21941 2748
rect 21965 2746 22021 2748
rect 21725 2694 21771 2746
rect 21771 2694 21781 2746
rect 21805 2694 21835 2746
rect 21835 2694 21847 2746
rect 21847 2694 21861 2746
rect 21885 2694 21899 2746
rect 21899 2694 21911 2746
rect 21911 2694 21941 2746
rect 21965 2694 21975 2746
rect 21975 2694 22021 2746
rect 21725 2692 21781 2694
rect 21805 2692 21861 2694
rect 21885 2692 21941 2694
rect 21965 2692 22021 2694
rect 22466 2488 22522 2544
rect 22282 2216 22338 2272
rect 23018 2352 23074 2408
rect 22190 1808 22246 1864
rect 21725 1658 21781 1660
rect 21805 1658 21861 1660
rect 21885 1658 21941 1660
rect 21965 1658 22021 1660
rect 21725 1606 21771 1658
rect 21771 1606 21781 1658
rect 21805 1606 21835 1658
rect 21835 1606 21847 1658
rect 21847 1606 21861 1658
rect 21885 1606 21899 1658
rect 21899 1606 21911 1658
rect 21911 1606 21941 1658
rect 21965 1606 21975 1658
rect 21975 1606 22021 1658
rect 21725 1604 21781 1606
rect 21805 1604 21861 1606
rect 21885 1604 21941 1606
rect 21965 1604 22021 1606
rect 24692 8730 24748 8732
rect 24772 8730 24828 8732
rect 24852 8730 24908 8732
rect 24932 8730 24988 8732
rect 24692 8678 24738 8730
rect 24738 8678 24748 8730
rect 24772 8678 24802 8730
rect 24802 8678 24814 8730
rect 24814 8678 24828 8730
rect 24852 8678 24866 8730
rect 24866 8678 24878 8730
rect 24878 8678 24908 8730
rect 24932 8678 24942 8730
rect 24942 8678 24988 8730
rect 24692 8676 24748 8678
rect 24772 8676 24828 8678
rect 24852 8676 24908 8678
rect 24932 8676 24988 8678
rect 24692 7642 24748 7644
rect 24772 7642 24828 7644
rect 24852 7642 24908 7644
rect 24932 7642 24988 7644
rect 24692 7590 24738 7642
rect 24738 7590 24748 7642
rect 24772 7590 24802 7642
rect 24802 7590 24814 7642
rect 24814 7590 24828 7642
rect 24852 7590 24866 7642
rect 24866 7590 24878 7642
rect 24878 7590 24908 7642
rect 24932 7590 24942 7642
rect 24942 7590 24988 7642
rect 24692 7588 24748 7590
rect 24772 7588 24828 7590
rect 24852 7588 24908 7590
rect 24932 7588 24988 7590
rect 24692 6554 24748 6556
rect 24772 6554 24828 6556
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 24692 6502 24738 6554
rect 24738 6502 24748 6554
rect 24772 6502 24802 6554
rect 24802 6502 24814 6554
rect 24814 6502 24828 6554
rect 24852 6502 24866 6554
rect 24866 6502 24878 6554
rect 24878 6502 24908 6554
rect 24932 6502 24942 6554
rect 24942 6502 24988 6554
rect 24692 6500 24748 6502
rect 24772 6500 24828 6502
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 24692 5466 24748 5468
rect 24772 5466 24828 5468
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 24692 5414 24738 5466
rect 24738 5414 24748 5466
rect 24772 5414 24802 5466
rect 24802 5414 24814 5466
rect 24814 5414 24828 5466
rect 24852 5414 24866 5466
rect 24866 5414 24878 5466
rect 24878 5414 24908 5466
rect 24932 5414 24942 5466
rect 24942 5414 24988 5466
rect 24692 5412 24748 5414
rect 24772 5412 24828 5414
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 24692 4378 24748 4380
rect 24772 4378 24828 4380
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 24692 4326 24738 4378
rect 24738 4326 24748 4378
rect 24772 4326 24802 4378
rect 24802 4326 24814 4378
rect 24814 4326 24828 4378
rect 24852 4326 24866 4378
rect 24866 4326 24878 4378
rect 24878 4326 24908 4378
rect 24932 4326 24942 4378
rect 24942 4326 24988 4378
rect 24692 4324 24748 4326
rect 24772 4324 24828 4326
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 24692 3290 24748 3292
rect 24772 3290 24828 3292
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 24692 3238 24738 3290
rect 24738 3238 24748 3290
rect 24772 3238 24802 3290
rect 24802 3238 24814 3290
rect 24814 3238 24828 3290
rect 24852 3238 24866 3290
rect 24866 3238 24878 3290
rect 24878 3238 24908 3290
rect 24932 3238 24942 3290
rect 24942 3238 24988 3290
rect 24692 3236 24748 3238
rect 24772 3236 24828 3238
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 24692 2202 24748 2204
rect 24772 2202 24828 2204
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 24692 2150 24738 2202
rect 24738 2150 24748 2202
rect 24772 2150 24802 2202
rect 24802 2150 24814 2202
rect 24814 2150 24828 2202
rect 24852 2150 24866 2202
rect 24866 2150 24878 2202
rect 24878 2150 24908 2202
rect 24932 2150 24942 2202
rect 24942 2150 24988 2202
rect 24692 2148 24748 2150
rect 24772 2148 24828 2150
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 24692 1114 24748 1116
rect 24772 1114 24828 1116
rect 24852 1114 24908 1116
rect 24932 1114 24988 1116
rect 24692 1062 24738 1114
rect 24738 1062 24748 1114
rect 24772 1062 24802 1114
rect 24802 1062 24814 1114
rect 24814 1062 24828 1114
rect 24852 1062 24866 1114
rect 24866 1062 24878 1114
rect 24878 1062 24908 1114
rect 24932 1062 24942 1114
rect 24942 1062 24988 1114
rect 24692 1060 24748 1062
rect 24772 1060 24828 1062
rect 24852 1060 24908 1062
rect 24932 1060 24988 1062
<< metal3 >>
rect 9765 9482 9831 9485
rect 11697 9482 11763 9485
rect 9765 9480 11763 9482
rect 9765 9424 9770 9480
rect 9826 9424 11702 9480
rect 11758 9424 11763 9480
rect 9765 9422 11763 9424
rect 9765 9419 9831 9422
rect 11697 9419 11763 9422
rect 6880 8736 7196 8737
rect 6880 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7196 8736
rect 6880 8671 7196 8672
rect 12814 8736 13130 8737
rect 12814 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13130 8736
rect 12814 8671 13130 8672
rect 18748 8736 19064 8737
rect 18748 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19064 8736
rect 18748 8671 19064 8672
rect 24682 8736 24998 8737
rect 24682 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 24998 8736
rect 24682 8671 24998 8672
rect 17861 8530 17927 8533
rect 18965 8530 19031 8533
rect 17861 8528 19031 8530
rect 17861 8472 17866 8528
rect 17922 8472 18970 8528
rect 19026 8472 19031 8528
rect 17861 8470 19031 8472
rect 17861 8467 17927 8470
rect 18965 8467 19031 8470
rect 10041 8394 10107 8397
rect 12985 8394 13051 8397
rect 10041 8392 13051 8394
rect 10041 8336 10046 8392
rect 10102 8336 12990 8392
rect 13046 8336 13051 8392
rect 10041 8334 13051 8336
rect 10041 8331 10107 8334
rect 12985 8331 13051 8334
rect 3913 8192 4229 8193
rect 3913 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4229 8192
rect 3913 8127 4229 8128
rect 9847 8192 10163 8193
rect 9847 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10163 8192
rect 9847 8127 10163 8128
rect 15781 8192 16097 8193
rect 15781 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16097 8192
rect 15781 8127 16097 8128
rect 21715 8192 22031 8193
rect 21715 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22031 8192
rect 21715 8127 22031 8128
rect 1945 7850 2011 7853
rect 15469 7850 15535 7853
rect 1945 7848 15535 7850
rect 1945 7792 1950 7848
rect 2006 7792 15474 7848
rect 15530 7792 15535 7848
rect 1945 7790 15535 7792
rect 1945 7787 2011 7790
rect 15469 7787 15535 7790
rect 6880 7648 7196 7649
rect 6880 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7196 7648
rect 6880 7583 7196 7584
rect 12814 7648 13130 7649
rect 12814 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13130 7648
rect 12814 7583 13130 7584
rect 18748 7648 19064 7649
rect 18748 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19064 7648
rect 18748 7583 19064 7584
rect 24682 7648 24998 7649
rect 24682 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 24998 7648
rect 24682 7583 24998 7584
rect 7373 7578 7439 7581
rect 10041 7578 10107 7581
rect 7373 7576 10107 7578
rect 7373 7520 7378 7576
rect 7434 7520 10046 7576
rect 10102 7520 10107 7576
rect 7373 7518 10107 7520
rect 7373 7515 7439 7518
rect 10041 7515 10107 7518
rect 5901 7442 5967 7445
rect 20069 7442 20135 7445
rect 5901 7440 20135 7442
rect 5901 7384 5906 7440
rect 5962 7384 20074 7440
rect 20130 7384 20135 7440
rect 5901 7382 20135 7384
rect 5901 7379 5967 7382
rect 20069 7379 20135 7382
rect 6177 7306 6243 7309
rect 19517 7306 19583 7309
rect 6177 7304 19583 7306
rect 6177 7248 6182 7304
rect 6238 7248 19522 7304
rect 19578 7248 19583 7304
rect 6177 7246 19583 7248
rect 6177 7243 6243 7246
rect 19517 7243 19583 7246
rect 3913 7104 4229 7105
rect 3913 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4229 7104
rect 3913 7039 4229 7040
rect 9847 7104 10163 7105
rect 9847 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10163 7104
rect 9847 7039 10163 7040
rect 15781 7104 16097 7105
rect 15781 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16097 7104
rect 15781 7039 16097 7040
rect 21715 7104 22031 7105
rect 21715 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22031 7104
rect 21715 7039 22031 7040
rect 6880 6560 7196 6561
rect 6880 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7196 6560
rect 6880 6495 7196 6496
rect 12814 6560 13130 6561
rect 12814 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13130 6560
rect 12814 6495 13130 6496
rect 18748 6560 19064 6561
rect 18748 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19064 6560
rect 18748 6495 19064 6496
rect 24682 6560 24998 6561
rect 24682 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 24998 6560
rect 24682 6495 24998 6496
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 9847 6016 10163 6017
rect 9847 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10163 6016
rect 9847 5951 10163 5952
rect 15781 6016 16097 6017
rect 15781 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16097 6016
rect 15781 5951 16097 5952
rect 21715 6016 22031 6017
rect 21715 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22031 6016
rect 21715 5951 22031 5952
rect 6880 5472 7196 5473
rect 6880 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7196 5472
rect 6880 5407 7196 5408
rect 12814 5472 13130 5473
rect 12814 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13130 5472
rect 12814 5407 13130 5408
rect 18748 5472 19064 5473
rect 18748 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19064 5472
rect 18748 5407 19064 5408
rect 24682 5472 24998 5473
rect 24682 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 24998 5472
rect 24682 5407 24998 5408
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 9847 4928 10163 4929
rect 9847 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10163 4928
rect 9847 4863 10163 4864
rect 15781 4928 16097 4929
rect 15781 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16097 4928
rect 15781 4863 16097 4864
rect 21715 4928 22031 4929
rect 21715 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22031 4928
rect 21715 4863 22031 4864
rect 6880 4384 7196 4385
rect 6880 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7196 4384
rect 6880 4319 7196 4320
rect 12814 4384 13130 4385
rect 12814 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13130 4384
rect 12814 4319 13130 4320
rect 18748 4384 19064 4385
rect 18748 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19064 4384
rect 18748 4319 19064 4320
rect 24682 4384 24998 4385
rect 24682 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 24998 4384
rect 24682 4319 24998 4320
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 9847 3840 10163 3841
rect 9847 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10163 3840
rect 9847 3775 10163 3776
rect 15781 3840 16097 3841
rect 15781 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16097 3840
rect 15781 3775 16097 3776
rect 21715 3840 22031 3841
rect 21715 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22031 3840
rect 21715 3775 22031 3776
rect 6880 3296 7196 3297
rect 6880 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7196 3296
rect 6880 3231 7196 3232
rect 12814 3296 13130 3297
rect 12814 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13130 3296
rect 12814 3231 13130 3232
rect 18748 3296 19064 3297
rect 18748 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19064 3296
rect 18748 3231 19064 3232
rect 24682 3296 24998 3297
rect 24682 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 24998 3296
rect 24682 3231 24998 3232
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 9847 2752 10163 2753
rect 9847 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10163 2752
rect 9847 2687 10163 2688
rect 15781 2752 16097 2753
rect 15781 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16097 2752
rect 15781 2687 16097 2688
rect 21715 2752 22031 2753
rect 21715 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22031 2752
rect 21715 2687 22031 2688
rect 11697 2546 11763 2549
rect 22461 2546 22527 2549
rect 11697 2544 22527 2546
rect 11697 2488 11702 2544
rect 11758 2488 22466 2544
rect 22522 2488 22527 2544
rect 11697 2486 22527 2488
rect 11697 2483 11763 2486
rect 22461 2483 22527 2486
rect 10225 2410 10291 2413
rect 23013 2410 23079 2413
rect 10225 2408 23079 2410
rect 10225 2352 10230 2408
rect 10286 2352 23018 2408
rect 23074 2352 23079 2408
rect 10225 2350 23079 2352
rect 10225 2347 10291 2350
rect 23013 2347 23079 2350
rect 22277 2274 22343 2277
rect 22050 2272 22343 2274
rect 22050 2216 22282 2272
rect 22338 2216 22343 2272
rect 22050 2214 22343 2216
rect 6880 2208 7196 2209
rect 6880 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7196 2208
rect 6880 2143 7196 2144
rect 12814 2208 13130 2209
rect 12814 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13130 2208
rect 12814 2143 13130 2144
rect 18748 2208 19064 2209
rect 18748 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19064 2208
rect 18748 2143 19064 2144
rect 9121 2002 9187 2005
rect 22050 2002 22110 2214
rect 22277 2211 22343 2214
rect 24682 2208 24998 2209
rect 24682 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 24998 2208
rect 24682 2143 24998 2144
rect 9121 2000 22110 2002
rect 9121 1944 9126 2000
rect 9182 1944 22110 2000
rect 9121 1942 22110 1944
rect 9121 1939 9187 1942
rect 7925 1866 7991 1869
rect 22185 1866 22251 1869
rect 7925 1864 22251 1866
rect 7925 1808 7930 1864
rect 7986 1808 22190 1864
rect 22246 1808 22251 1864
rect 7925 1806 22251 1808
rect 7925 1803 7991 1806
rect 22185 1803 22251 1806
rect 3913 1664 4229 1665
rect 3913 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4229 1664
rect 3913 1599 4229 1600
rect 9847 1664 10163 1665
rect 9847 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10163 1664
rect 9847 1599 10163 1600
rect 15781 1664 16097 1665
rect 15781 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16097 1664
rect 15781 1599 16097 1600
rect 21715 1664 22031 1665
rect 21715 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22031 1664
rect 21715 1599 22031 1600
rect 6880 1120 7196 1121
rect 6880 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7196 1120
rect 6880 1055 7196 1056
rect 12814 1120 13130 1121
rect 12814 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13130 1120
rect 12814 1055 13130 1056
rect 18748 1120 19064 1121
rect 18748 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19064 1120
rect 18748 1055 19064 1056
rect 24682 1120 24998 1121
rect 24682 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 24998 1120
rect 24682 1055 24998 1056
<< via3 >>
rect 6886 8732 6950 8736
rect 6886 8676 6890 8732
rect 6890 8676 6946 8732
rect 6946 8676 6950 8732
rect 6886 8672 6950 8676
rect 6966 8732 7030 8736
rect 6966 8676 6970 8732
rect 6970 8676 7026 8732
rect 7026 8676 7030 8732
rect 6966 8672 7030 8676
rect 7046 8732 7110 8736
rect 7046 8676 7050 8732
rect 7050 8676 7106 8732
rect 7106 8676 7110 8732
rect 7046 8672 7110 8676
rect 7126 8732 7190 8736
rect 7126 8676 7130 8732
rect 7130 8676 7186 8732
rect 7186 8676 7190 8732
rect 7126 8672 7190 8676
rect 12820 8732 12884 8736
rect 12820 8676 12824 8732
rect 12824 8676 12880 8732
rect 12880 8676 12884 8732
rect 12820 8672 12884 8676
rect 12900 8732 12964 8736
rect 12900 8676 12904 8732
rect 12904 8676 12960 8732
rect 12960 8676 12964 8732
rect 12900 8672 12964 8676
rect 12980 8732 13044 8736
rect 12980 8676 12984 8732
rect 12984 8676 13040 8732
rect 13040 8676 13044 8732
rect 12980 8672 13044 8676
rect 13060 8732 13124 8736
rect 13060 8676 13064 8732
rect 13064 8676 13120 8732
rect 13120 8676 13124 8732
rect 13060 8672 13124 8676
rect 18754 8732 18818 8736
rect 18754 8676 18758 8732
rect 18758 8676 18814 8732
rect 18814 8676 18818 8732
rect 18754 8672 18818 8676
rect 18834 8732 18898 8736
rect 18834 8676 18838 8732
rect 18838 8676 18894 8732
rect 18894 8676 18898 8732
rect 18834 8672 18898 8676
rect 18914 8732 18978 8736
rect 18914 8676 18918 8732
rect 18918 8676 18974 8732
rect 18974 8676 18978 8732
rect 18914 8672 18978 8676
rect 18994 8732 19058 8736
rect 18994 8676 18998 8732
rect 18998 8676 19054 8732
rect 19054 8676 19058 8732
rect 18994 8672 19058 8676
rect 24688 8732 24752 8736
rect 24688 8676 24692 8732
rect 24692 8676 24748 8732
rect 24748 8676 24752 8732
rect 24688 8672 24752 8676
rect 24768 8732 24832 8736
rect 24768 8676 24772 8732
rect 24772 8676 24828 8732
rect 24828 8676 24832 8732
rect 24768 8672 24832 8676
rect 24848 8732 24912 8736
rect 24848 8676 24852 8732
rect 24852 8676 24908 8732
rect 24908 8676 24912 8732
rect 24848 8672 24912 8676
rect 24928 8732 24992 8736
rect 24928 8676 24932 8732
rect 24932 8676 24988 8732
rect 24988 8676 24992 8732
rect 24928 8672 24992 8676
rect 3919 8188 3983 8192
rect 3919 8132 3923 8188
rect 3923 8132 3979 8188
rect 3979 8132 3983 8188
rect 3919 8128 3983 8132
rect 3999 8188 4063 8192
rect 3999 8132 4003 8188
rect 4003 8132 4059 8188
rect 4059 8132 4063 8188
rect 3999 8128 4063 8132
rect 4079 8188 4143 8192
rect 4079 8132 4083 8188
rect 4083 8132 4139 8188
rect 4139 8132 4143 8188
rect 4079 8128 4143 8132
rect 4159 8188 4223 8192
rect 4159 8132 4163 8188
rect 4163 8132 4219 8188
rect 4219 8132 4223 8188
rect 4159 8128 4223 8132
rect 9853 8188 9917 8192
rect 9853 8132 9857 8188
rect 9857 8132 9913 8188
rect 9913 8132 9917 8188
rect 9853 8128 9917 8132
rect 9933 8188 9997 8192
rect 9933 8132 9937 8188
rect 9937 8132 9993 8188
rect 9993 8132 9997 8188
rect 9933 8128 9997 8132
rect 10013 8188 10077 8192
rect 10013 8132 10017 8188
rect 10017 8132 10073 8188
rect 10073 8132 10077 8188
rect 10013 8128 10077 8132
rect 10093 8188 10157 8192
rect 10093 8132 10097 8188
rect 10097 8132 10153 8188
rect 10153 8132 10157 8188
rect 10093 8128 10157 8132
rect 15787 8188 15851 8192
rect 15787 8132 15791 8188
rect 15791 8132 15847 8188
rect 15847 8132 15851 8188
rect 15787 8128 15851 8132
rect 15867 8188 15931 8192
rect 15867 8132 15871 8188
rect 15871 8132 15927 8188
rect 15927 8132 15931 8188
rect 15867 8128 15931 8132
rect 15947 8188 16011 8192
rect 15947 8132 15951 8188
rect 15951 8132 16007 8188
rect 16007 8132 16011 8188
rect 15947 8128 16011 8132
rect 16027 8188 16091 8192
rect 16027 8132 16031 8188
rect 16031 8132 16087 8188
rect 16087 8132 16091 8188
rect 16027 8128 16091 8132
rect 21721 8188 21785 8192
rect 21721 8132 21725 8188
rect 21725 8132 21781 8188
rect 21781 8132 21785 8188
rect 21721 8128 21785 8132
rect 21801 8188 21865 8192
rect 21801 8132 21805 8188
rect 21805 8132 21861 8188
rect 21861 8132 21865 8188
rect 21801 8128 21865 8132
rect 21881 8188 21945 8192
rect 21881 8132 21885 8188
rect 21885 8132 21941 8188
rect 21941 8132 21945 8188
rect 21881 8128 21945 8132
rect 21961 8188 22025 8192
rect 21961 8132 21965 8188
rect 21965 8132 22021 8188
rect 22021 8132 22025 8188
rect 21961 8128 22025 8132
rect 6886 7644 6950 7648
rect 6886 7588 6890 7644
rect 6890 7588 6946 7644
rect 6946 7588 6950 7644
rect 6886 7584 6950 7588
rect 6966 7644 7030 7648
rect 6966 7588 6970 7644
rect 6970 7588 7026 7644
rect 7026 7588 7030 7644
rect 6966 7584 7030 7588
rect 7046 7644 7110 7648
rect 7046 7588 7050 7644
rect 7050 7588 7106 7644
rect 7106 7588 7110 7644
rect 7046 7584 7110 7588
rect 7126 7644 7190 7648
rect 7126 7588 7130 7644
rect 7130 7588 7186 7644
rect 7186 7588 7190 7644
rect 7126 7584 7190 7588
rect 12820 7644 12884 7648
rect 12820 7588 12824 7644
rect 12824 7588 12880 7644
rect 12880 7588 12884 7644
rect 12820 7584 12884 7588
rect 12900 7644 12964 7648
rect 12900 7588 12904 7644
rect 12904 7588 12960 7644
rect 12960 7588 12964 7644
rect 12900 7584 12964 7588
rect 12980 7644 13044 7648
rect 12980 7588 12984 7644
rect 12984 7588 13040 7644
rect 13040 7588 13044 7644
rect 12980 7584 13044 7588
rect 13060 7644 13124 7648
rect 13060 7588 13064 7644
rect 13064 7588 13120 7644
rect 13120 7588 13124 7644
rect 13060 7584 13124 7588
rect 18754 7644 18818 7648
rect 18754 7588 18758 7644
rect 18758 7588 18814 7644
rect 18814 7588 18818 7644
rect 18754 7584 18818 7588
rect 18834 7644 18898 7648
rect 18834 7588 18838 7644
rect 18838 7588 18894 7644
rect 18894 7588 18898 7644
rect 18834 7584 18898 7588
rect 18914 7644 18978 7648
rect 18914 7588 18918 7644
rect 18918 7588 18974 7644
rect 18974 7588 18978 7644
rect 18914 7584 18978 7588
rect 18994 7644 19058 7648
rect 18994 7588 18998 7644
rect 18998 7588 19054 7644
rect 19054 7588 19058 7644
rect 18994 7584 19058 7588
rect 24688 7644 24752 7648
rect 24688 7588 24692 7644
rect 24692 7588 24748 7644
rect 24748 7588 24752 7644
rect 24688 7584 24752 7588
rect 24768 7644 24832 7648
rect 24768 7588 24772 7644
rect 24772 7588 24828 7644
rect 24828 7588 24832 7644
rect 24768 7584 24832 7588
rect 24848 7644 24912 7648
rect 24848 7588 24852 7644
rect 24852 7588 24908 7644
rect 24908 7588 24912 7644
rect 24848 7584 24912 7588
rect 24928 7644 24992 7648
rect 24928 7588 24932 7644
rect 24932 7588 24988 7644
rect 24988 7588 24992 7644
rect 24928 7584 24992 7588
rect 3919 7100 3983 7104
rect 3919 7044 3923 7100
rect 3923 7044 3979 7100
rect 3979 7044 3983 7100
rect 3919 7040 3983 7044
rect 3999 7100 4063 7104
rect 3999 7044 4003 7100
rect 4003 7044 4059 7100
rect 4059 7044 4063 7100
rect 3999 7040 4063 7044
rect 4079 7100 4143 7104
rect 4079 7044 4083 7100
rect 4083 7044 4139 7100
rect 4139 7044 4143 7100
rect 4079 7040 4143 7044
rect 4159 7100 4223 7104
rect 4159 7044 4163 7100
rect 4163 7044 4219 7100
rect 4219 7044 4223 7100
rect 4159 7040 4223 7044
rect 9853 7100 9917 7104
rect 9853 7044 9857 7100
rect 9857 7044 9913 7100
rect 9913 7044 9917 7100
rect 9853 7040 9917 7044
rect 9933 7100 9997 7104
rect 9933 7044 9937 7100
rect 9937 7044 9993 7100
rect 9993 7044 9997 7100
rect 9933 7040 9997 7044
rect 10013 7100 10077 7104
rect 10013 7044 10017 7100
rect 10017 7044 10073 7100
rect 10073 7044 10077 7100
rect 10013 7040 10077 7044
rect 10093 7100 10157 7104
rect 10093 7044 10097 7100
rect 10097 7044 10153 7100
rect 10153 7044 10157 7100
rect 10093 7040 10157 7044
rect 15787 7100 15851 7104
rect 15787 7044 15791 7100
rect 15791 7044 15847 7100
rect 15847 7044 15851 7100
rect 15787 7040 15851 7044
rect 15867 7100 15931 7104
rect 15867 7044 15871 7100
rect 15871 7044 15927 7100
rect 15927 7044 15931 7100
rect 15867 7040 15931 7044
rect 15947 7100 16011 7104
rect 15947 7044 15951 7100
rect 15951 7044 16007 7100
rect 16007 7044 16011 7100
rect 15947 7040 16011 7044
rect 16027 7100 16091 7104
rect 16027 7044 16031 7100
rect 16031 7044 16087 7100
rect 16087 7044 16091 7100
rect 16027 7040 16091 7044
rect 21721 7100 21785 7104
rect 21721 7044 21725 7100
rect 21725 7044 21781 7100
rect 21781 7044 21785 7100
rect 21721 7040 21785 7044
rect 21801 7100 21865 7104
rect 21801 7044 21805 7100
rect 21805 7044 21861 7100
rect 21861 7044 21865 7100
rect 21801 7040 21865 7044
rect 21881 7100 21945 7104
rect 21881 7044 21885 7100
rect 21885 7044 21941 7100
rect 21941 7044 21945 7100
rect 21881 7040 21945 7044
rect 21961 7100 22025 7104
rect 21961 7044 21965 7100
rect 21965 7044 22021 7100
rect 22021 7044 22025 7100
rect 21961 7040 22025 7044
rect 6886 6556 6950 6560
rect 6886 6500 6890 6556
rect 6890 6500 6946 6556
rect 6946 6500 6950 6556
rect 6886 6496 6950 6500
rect 6966 6556 7030 6560
rect 6966 6500 6970 6556
rect 6970 6500 7026 6556
rect 7026 6500 7030 6556
rect 6966 6496 7030 6500
rect 7046 6556 7110 6560
rect 7046 6500 7050 6556
rect 7050 6500 7106 6556
rect 7106 6500 7110 6556
rect 7046 6496 7110 6500
rect 7126 6556 7190 6560
rect 7126 6500 7130 6556
rect 7130 6500 7186 6556
rect 7186 6500 7190 6556
rect 7126 6496 7190 6500
rect 12820 6556 12884 6560
rect 12820 6500 12824 6556
rect 12824 6500 12880 6556
rect 12880 6500 12884 6556
rect 12820 6496 12884 6500
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 18754 6556 18818 6560
rect 18754 6500 18758 6556
rect 18758 6500 18814 6556
rect 18814 6500 18818 6556
rect 18754 6496 18818 6500
rect 18834 6556 18898 6560
rect 18834 6500 18838 6556
rect 18838 6500 18894 6556
rect 18894 6500 18898 6556
rect 18834 6496 18898 6500
rect 18914 6556 18978 6560
rect 18914 6500 18918 6556
rect 18918 6500 18974 6556
rect 18974 6500 18978 6556
rect 18914 6496 18978 6500
rect 18994 6556 19058 6560
rect 18994 6500 18998 6556
rect 18998 6500 19054 6556
rect 19054 6500 19058 6556
rect 18994 6496 19058 6500
rect 24688 6556 24752 6560
rect 24688 6500 24692 6556
rect 24692 6500 24748 6556
rect 24748 6500 24752 6556
rect 24688 6496 24752 6500
rect 24768 6556 24832 6560
rect 24768 6500 24772 6556
rect 24772 6500 24828 6556
rect 24828 6500 24832 6556
rect 24768 6496 24832 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 9853 6012 9917 6016
rect 9853 5956 9857 6012
rect 9857 5956 9913 6012
rect 9913 5956 9917 6012
rect 9853 5952 9917 5956
rect 9933 6012 9997 6016
rect 9933 5956 9937 6012
rect 9937 5956 9993 6012
rect 9993 5956 9997 6012
rect 9933 5952 9997 5956
rect 10013 6012 10077 6016
rect 10013 5956 10017 6012
rect 10017 5956 10073 6012
rect 10073 5956 10077 6012
rect 10013 5952 10077 5956
rect 10093 6012 10157 6016
rect 10093 5956 10097 6012
rect 10097 5956 10153 6012
rect 10153 5956 10157 6012
rect 10093 5952 10157 5956
rect 15787 6012 15851 6016
rect 15787 5956 15791 6012
rect 15791 5956 15847 6012
rect 15847 5956 15851 6012
rect 15787 5952 15851 5956
rect 15867 6012 15931 6016
rect 15867 5956 15871 6012
rect 15871 5956 15927 6012
rect 15927 5956 15931 6012
rect 15867 5952 15931 5956
rect 15947 6012 16011 6016
rect 15947 5956 15951 6012
rect 15951 5956 16007 6012
rect 16007 5956 16011 6012
rect 15947 5952 16011 5956
rect 16027 6012 16091 6016
rect 16027 5956 16031 6012
rect 16031 5956 16087 6012
rect 16087 5956 16091 6012
rect 16027 5952 16091 5956
rect 21721 6012 21785 6016
rect 21721 5956 21725 6012
rect 21725 5956 21781 6012
rect 21781 5956 21785 6012
rect 21721 5952 21785 5956
rect 21801 6012 21865 6016
rect 21801 5956 21805 6012
rect 21805 5956 21861 6012
rect 21861 5956 21865 6012
rect 21801 5952 21865 5956
rect 21881 6012 21945 6016
rect 21881 5956 21885 6012
rect 21885 5956 21941 6012
rect 21941 5956 21945 6012
rect 21881 5952 21945 5956
rect 21961 6012 22025 6016
rect 21961 5956 21965 6012
rect 21965 5956 22021 6012
rect 22021 5956 22025 6012
rect 21961 5952 22025 5956
rect 6886 5468 6950 5472
rect 6886 5412 6890 5468
rect 6890 5412 6946 5468
rect 6946 5412 6950 5468
rect 6886 5408 6950 5412
rect 6966 5468 7030 5472
rect 6966 5412 6970 5468
rect 6970 5412 7026 5468
rect 7026 5412 7030 5468
rect 6966 5408 7030 5412
rect 7046 5468 7110 5472
rect 7046 5412 7050 5468
rect 7050 5412 7106 5468
rect 7106 5412 7110 5468
rect 7046 5408 7110 5412
rect 7126 5468 7190 5472
rect 7126 5412 7130 5468
rect 7130 5412 7186 5468
rect 7186 5412 7190 5468
rect 7126 5408 7190 5412
rect 12820 5468 12884 5472
rect 12820 5412 12824 5468
rect 12824 5412 12880 5468
rect 12880 5412 12884 5468
rect 12820 5408 12884 5412
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 18754 5468 18818 5472
rect 18754 5412 18758 5468
rect 18758 5412 18814 5468
rect 18814 5412 18818 5468
rect 18754 5408 18818 5412
rect 18834 5468 18898 5472
rect 18834 5412 18838 5468
rect 18838 5412 18894 5468
rect 18894 5412 18898 5468
rect 18834 5408 18898 5412
rect 18914 5468 18978 5472
rect 18914 5412 18918 5468
rect 18918 5412 18974 5468
rect 18974 5412 18978 5468
rect 18914 5408 18978 5412
rect 18994 5468 19058 5472
rect 18994 5412 18998 5468
rect 18998 5412 19054 5468
rect 19054 5412 19058 5468
rect 18994 5408 19058 5412
rect 24688 5468 24752 5472
rect 24688 5412 24692 5468
rect 24692 5412 24748 5468
rect 24748 5412 24752 5468
rect 24688 5408 24752 5412
rect 24768 5468 24832 5472
rect 24768 5412 24772 5468
rect 24772 5412 24828 5468
rect 24828 5412 24832 5468
rect 24768 5408 24832 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 9853 4924 9917 4928
rect 9853 4868 9857 4924
rect 9857 4868 9913 4924
rect 9913 4868 9917 4924
rect 9853 4864 9917 4868
rect 9933 4924 9997 4928
rect 9933 4868 9937 4924
rect 9937 4868 9993 4924
rect 9993 4868 9997 4924
rect 9933 4864 9997 4868
rect 10013 4924 10077 4928
rect 10013 4868 10017 4924
rect 10017 4868 10073 4924
rect 10073 4868 10077 4924
rect 10013 4864 10077 4868
rect 10093 4924 10157 4928
rect 10093 4868 10097 4924
rect 10097 4868 10153 4924
rect 10153 4868 10157 4924
rect 10093 4864 10157 4868
rect 15787 4924 15851 4928
rect 15787 4868 15791 4924
rect 15791 4868 15847 4924
rect 15847 4868 15851 4924
rect 15787 4864 15851 4868
rect 15867 4924 15931 4928
rect 15867 4868 15871 4924
rect 15871 4868 15927 4924
rect 15927 4868 15931 4924
rect 15867 4864 15931 4868
rect 15947 4924 16011 4928
rect 15947 4868 15951 4924
rect 15951 4868 16007 4924
rect 16007 4868 16011 4924
rect 15947 4864 16011 4868
rect 16027 4924 16091 4928
rect 16027 4868 16031 4924
rect 16031 4868 16087 4924
rect 16087 4868 16091 4924
rect 16027 4864 16091 4868
rect 21721 4924 21785 4928
rect 21721 4868 21725 4924
rect 21725 4868 21781 4924
rect 21781 4868 21785 4924
rect 21721 4864 21785 4868
rect 21801 4924 21865 4928
rect 21801 4868 21805 4924
rect 21805 4868 21861 4924
rect 21861 4868 21865 4924
rect 21801 4864 21865 4868
rect 21881 4924 21945 4928
rect 21881 4868 21885 4924
rect 21885 4868 21941 4924
rect 21941 4868 21945 4924
rect 21881 4864 21945 4868
rect 21961 4924 22025 4928
rect 21961 4868 21965 4924
rect 21965 4868 22021 4924
rect 22021 4868 22025 4924
rect 21961 4864 22025 4868
rect 6886 4380 6950 4384
rect 6886 4324 6890 4380
rect 6890 4324 6946 4380
rect 6946 4324 6950 4380
rect 6886 4320 6950 4324
rect 6966 4380 7030 4384
rect 6966 4324 6970 4380
rect 6970 4324 7026 4380
rect 7026 4324 7030 4380
rect 6966 4320 7030 4324
rect 7046 4380 7110 4384
rect 7046 4324 7050 4380
rect 7050 4324 7106 4380
rect 7106 4324 7110 4380
rect 7046 4320 7110 4324
rect 7126 4380 7190 4384
rect 7126 4324 7130 4380
rect 7130 4324 7186 4380
rect 7186 4324 7190 4380
rect 7126 4320 7190 4324
rect 12820 4380 12884 4384
rect 12820 4324 12824 4380
rect 12824 4324 12880 4380
rect 12880 4324 12884 4380
rect 12820 4320 12884 4324
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 18754 4380 18818 4384
rect 18754 4324 18758 4380
rect 18758 4324 18814 4380
rect 18814 4324 18818 4380
rect 18754 4320 18818 4324
rect 18834 4380 18898 4384
rect 18834 4324 18838 4380
rect 18838 4324 18894 4380
rect 18894 4324 18898 4380
rect 18834 4320 18898 4324
rect 18914 4380 18978 4384
rect 18914 4324 18918 4380
rect 18918 4324 18974 4380
rect 18974 4324 18978 4380
rect 18914 4320 18978 4324
rect 18994 4380 19058 4384
rect 18994 4324 18998 4380
rect 18998 4324 19054 4380
rect 19054 4324 19058 4380
rect 18994 4320 19058 4324
rect 24688 4380 24752 4384
rect 24688 4324 24692 4380
rect 24692 4324 24748 4380
rect 24748 4324 24752 4380
rect 24688 4320 24752 4324
rect 24768 4380 24832 4384
rect 24768 4324 24772 4380
rect 24772 4324 24828 4380
rect 24828 4324 24832 4380
rect 24768 4320 24832 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 9853 3836 9917 3840
rect 9853 3780 9857 3836
rect 9857 3780 9913 3836
rect 9913 3780 9917 3836
rect 9853 3776 9917 3780
rect 9933 3836 9997 3840
rect 9933 3780 9937 3836
rect 9937 3780 9993 3836
rect 9993 3780 9997 3836
rect 9933 3776 9997 3780
rect 10013 3836 10077 3840
rect 10013 3780 10017 3836
rect 10017 3780 10073 3836
rect 10073 3780 10077 3836
rect 10013 3776 10077 3780
rect 10093 3836 10157 3840
rect 10093 3780 10097 3836
rect 10097 3780 10153 3836
rect 10153 3780 10157 3836
rect 10093 3776 10157 3780
rect 15787 3836 15851 3840
rect 15787 3780 15791 3836
rect 15791 3780 15847 3836
rect 15847 3780 15851 3836
rect 15787 3776 15851 3780
rect 15867 3836 15931 3840
rect 15867 3780 15871 3836
rect 15871 3780 15927 3836
rect 15927 3780 15931 3836
rect 15867 3776 15931 3780
rect 15947 3836 16011 3840
rect 15947 3780 15951 3836
rect 15951 3780 16007 3836
rect 16007 3780 16011 3836
rect 15947 3776 16011 3780
rect 16027 3836 16091 3840
rect 16027 3780 16031 3836
rect 16031 3780 16087 3836
rect 16087 3780 16091 3836
rect 16027 3776 16091 3780
rect 21721 3836 21785 3840
rect 21721 3780 21725 3836
rect 21725 3780 21781 3836
rect 21781 3780 21785 3836
rect 21721 3776 21785 3780
rect 21801 3836 21865 3840
rect 21801 3780 21805 3836
rect 21805 3780 21861 3836
rect 21861 3780 21865 3836
rect 21801 3776 21865 3780
rect 21881 3836 21945 3840
rect 21881 3780 21885 3836
rect 21885 3780 21941 3836
rect 21941 3780 21945 3836
rect 21881 3776 21945 3780
rect 21961 3836 22025 3840
rect 21961 3780 21965 3836
rect 21965 3780 22021 3836
rect 22021 3780 22025 3836
rect 21961 3776 22025 3780
rect 6886 3292 6950 3296
rect 6886 3236 6890 3292
rect 6890 3236 6946 3292
rect 6946 3236 6950 3292
rect 6886 3232 6950 3236
rect 6966 3292 7030 3296
rect 6966 3236 6970 3292
rect 6970 3236 7026 3292
rect 7026 3236 7030 3292
rect 6966 3232 7030 3236
rect 7046 3292 7110 3296
rect 7046 3236 7050 3292
rect 7050 3236 7106 3292
rect 7106 3236 7110 3292
rect 7046 3232 7110 3236
rect 7126 3292 7190 3296
rect 7126 3236 7130 3292
rect 7130 3236 7186 3292
rect 7186 3236 7190 3292
rect 7126 3232 7190 3236
rect 12820 3292 12884 3296
rect 12820 3236 12824 3292
rect 12824 3236 12880 3292
rect 12880 3236 12884 3292
rect 12820 3232 12884 3236
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 18754 3292 18818 3296
rect 18754 3236 18758 3292
rect 18758 3236 18814 3292
rect 18814 3236 18818 3292
rect 18754 3232 18818 3236
rect 18834 3292 18898 3296
rect 18834 3236 18838 3292
rect 18838 3236 18894 3292
rect 18894 3236 18898 3292
rect 18834 3232 18898 3236
rect 18914 3292 18978 3296
rect 18914 3236 18918 3292
rect 18918 3236 18974 3292
rect 18974 3236 18978 3292
rect 18914 3232 18978 3236
rect 18994 3292 19058 3296
rect 18994 3236 18998 3292
rect 18998 3236 19054 3292
rect 19054 3236 19058 3292
rect 18994 3232 19058 3236
rect 24688 3292 24752 3296
rect 24688 3236 24692 3292
rect 24692 3236 24748 3292
rect 24748 3236 24752 3292
rect 24688 3232 24752 3236
rect 24768 3292 24832 3296
rect 24768 3236 24772 3292
rect 24772 3236 24828 3292
rect 24828 3236 24832 3292
rect 24768 3232 24832 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 9853 2748 9917 2752
rect 9853 2692 9857 2748
rect 9857 2692 9913 2748
rect 9913 2692 9917 2748
rect 9853 2688 9917 2692
rect 9933 2748 9997 2752
rect 9933 2692 9937 2748
rect 9937 2692 9993 2748
rect 9993 2692 9997 2748
rect 9933 2688 9997 2692
rect 10013 2748 10077 2752
rect 10013 2692 10017 2748
rect 10017 2692 10073 2748
rect 10073 2692 10077 2748
rect 10013 2688 10077 2692
rect 10093 2748 10157 2752
rect 10093 2692 10097 2748
rect 10097 2692 10153 2748
rect 10153 2692 10157 2748
rect 10093 2688 10157 2692
rect 15787 2748 15851 2752
rect 15787 2692 15791 2748
rect 15791 2692 15847 2748
rect 15847 2692 15851 2748
rect 15787 2688 15851 2692
rect 15867 2748 15931 2752
rect 15867 2692 15871 2748
rect 15871 2692 15927 2748
rect 15927 2692 15931 2748
rect 15867 2688 15931 2692
rect 15947 2748 16011 2752
rect 15947 2692 15951 2748
rect 15951 2692 16007 2748
rect 16007 2692 16011 2748
rect 15947 2688 16011 2692
rect 16027 2748 16091 2752
rect 16027 2692 16031 2748
rect 16031 2692 16087 2748
rect 16087 2692 16091 2748
rect 16027 2688 16091 2692
rect 21721 2748 21785 2752
rect 21721 2692 21725 2748
rect 21725 2692 21781 2748
rect 21781 2692 21785 2748
rect 21721 2688 21785 2692
rect 21801 2748 21865 2752
rect 21801 2692 21805 2748
rect 21805 2692 21861 2748
rect 21861 2692 21865 2748
rect 21801 2688 21865 2692
rect 21881 2748 21945 2752
rect 21881 2692 21885 2748
rect 21885 2692 21941 2748
rect 21941 2692 21945 2748
rect 21881 2688 21945 2692
rect 21961 2748 22025 2752
rect 21961 2692 21965 2748
rect 21965 2692 22021 2748
rect 22021 2692 22025 2748
rect 21961 2688 22025 2692
rect 6886 2204 6950 2208
rect 6886 2148 6890 2204
rect 6890 2148 6946 2204
rect 6946 2148 6950 2204
rect 6886 2144 6950 2148
rect 6966 2204 7030 2208
rect 6966 2148 6970 2204
rect 6970 2148 7026 2204
rect 7026 2148 7030 2204
rect 6966 2144 7030 2148
rect 7046 2204 7110 2208
rect 7046 2148 7050 2204
rect 7050 2148 7106 2204
rect 7106 2148 7110 2204
rect 7046 2144 7110 2148
rect 7126 2204 7190 2208
rect 7126 2148 7130 2204
rect 7130 2148 7186 2204
rect 7186 2148 7190 2204
rect 7126 2144 7190 2148
rect 12820 2204 12884 2208
rect 12820 2148 12824 2204
rect 12824 2148 12880 2204
rect 12880 2148 12884 2204
rect 12820 2144 12884 2148
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 18754 2204 18818 2208
rect 18754 2148 18758 2204
rect 18758 2148 18814 2204
rect 18814 2148 18818 2204
rect 18754 2144 18818 2148
rect 18834 2204 18898 2208
rect 18834 2148 18838 2204
rect 18838 2148 18894 2204
rect 18894 2148 18898 2204
rect 18834 2144 18898 2148
rect 18914 2204 18978 2208
rect 18914 2148 18918 2204
rect 18918 2148 18974 2204
rect 18974 2148 18978 2204
rect 18914 2144 18978 2148
rect 18994 2204 19058 2208
rect 18994 2148 18998 2204
rect 18998 2148 19054 2204
rect 19054 2148 19058 2204
rect 18994 2144 19058 2148
rect 24688 2204 24752 2208
rect 24688 2148 24692 2204
rect 24692 2148 24748 2204
rect 24748 2148 24752 2204
rect 24688 2144 24752 2148
rect 24768 2204 24832 2208
rect 24768 2148 24772 2204
rect 24772 2148 24828 2204
rect 24828 2148 24832 2204
rect 24768 2144 24832 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 3919 1660 3983 1664
rect 3919 1604 3923 1660
rect 3923 1604 3979 1660
rect 3979 1604 3983 1660
rect 3919 1600 3983 1604
rect 3999 1660 4063 1664
rect 3999 1604 4003 1660
rect 4003 1604 4059 1660
rect 4059 1604 4063 1660
rect 3999 1600 4063 1604
rect 4079 1660 4143 1664
rect 4079 1604 4083 1660
rect 4083 1604 4139 1660
rect 4139 1604 4143 1660
rect 4079 1600 4143 1604
rect 4159 1660 4223 1664
rect 4159 1604 4163 1660
rect 4163 1604 4219 1660
rect 4219 1604 4223 1660
rect 4159 1600 4223 1604
rect 9853 1660 9917 1664
rect 9853 1604 9857 1660
rect 9857 1604 9913 1660
rect 9913 1604 9917 1660
rect 9853 1600 9917 1604
rect 9933 1660 9997 1664
rect 9933 1604 9937 1660
rect 9937 1604 9993 1660
rect 9993 1604 9997 1660
rect 9933 1600 9997 1604
rect 10013 1660 10077 1664
rect 10013 1604 10017 1660
rect 10017 1604 10073 1660
rect 10073 1604 10077 1660
rect 10013 1600 10077 1604
rect 10093 1660 10157 1664
rect 10093 1604 10097 1660
rect 10097 1604 10153 1660
rect 10153 1604 10157 1660
rect 10093 1600 10157 1604
rect 15787 1660 15851 1664
rect 15787 1604 15791 1660
rect 15791 1604 15847 1660
rect 15847 1604 15851 1660
rect 15787 1600 15851 1604
rect 15867 1660 15931 1664
rect 15867 1604 15871 1660
rect 15871 1604 15927 1660
rect 15927 1604 15931 1660
rect 15867 1600 15931 1604
rect 15947 1660 16011 1664
rect 15947 1604 15951 1660
rect 15951 1604 16007 1660
rect 16007 1604 16011 1660
rect 15947 1600 16011 1604
rect 16027 1660 16091 1664
rect 16027 1604 16031 1660
rect 16031 1604 16087 1660
rect 16087 1604 16091 1660
rect 16027 1600 16091 1604
rect 21721 1660 21785 1664
rect 21721 1604 21725 1660
rect 21725 1604 21781 1660
rect 21781 1604 21785 1660
rect 21721 1600 21785 1604
rect 21801 1660 21865 1664
rect 21801 1604 21805 1660
rect 21805 1604 21861 1660
rect 21861 1604 21865 1660
rect 21801 1600 21865 1604
rect 21881 1660 21945 1664
rect 21881 1604 21885 1660
rect 21885 1604 21941 1660
rect 21941 1604 21945 1660
rect 21881 1600 21945 1604
rect 21961 1660 22025 1664
rect 21961 1604 21965 1660
rect 21965 1604 22021 1660
rect 22021 1604 22025 1660
rect 21961 1600 22025 1604
rect 6886 1116 6950 1120
rect 6886 1060 6890 1116
rect 6890 1060 6946 1116
rect 6946 1060 6950 1116
rect 6886 1056 6950 1060
rect 6966 1116 7030 1120
rect 6966 1060 6970 1116
rect 6970 1060 7026 1116
rect 7026 1060 7030 1116
rect 6966 1056 7030 1060
rect 7046 1116 7110 1120
rect 7046 1060 7050 1116
rect 7050 1060 7106 1116
rect 7106 1060 7110 1116
rect 7046 1056 7110 1060
rect 7126 1116 7190 1120
rect 7126 1060 7130 1116
rect 7130 1060 7186 1116
rect 7186 1060 7190 1116
rect 7126 1056 7190 1060
rect 12820 1116 12884 1120
rect 12820 1060 12824 1116
rect 12824 1060 12880 1116
rect 12880 1060 12884 1116
rect 12820 1056 12884 1060
rect 12900 1116 12964 1120
rect 12900 1060 12904 1116
rect 12904 1060 12960 1116
rect 12960 1060 12964 1116
rect 12900 1056 12964 1060
rect 12980 1116 13044 1120
rect 12980 1060 12984 1116
rect 12984 1060 13040 1116
rect 13040 1060 13044 1116
rect 12980 1056 13044 1060
rect 13060 1116 13124 1120
rect 13060 1060 13064 1116
rect 13064 1060 13120 1116
rect 13120 1060 13124 1116
rect 13060 1056 13124 1060
rect 18754 1116 18818 1120
rect 18754 1060 18758 1116
rect 18758 1060 18814 1116
rect 18814 1060 18818 1116
rect 18754 1056 18818 1060
rect 18834 1116 18898 1120
rect 18834 1060 18838 1116
rect 18838 1060 18894 1116
rect 18894 1060 18898 1116
rect 18834 1056 18898 1060
rect 18914 1116 18978 1120
rect 18914 1060 18918 1116
rect 18918 1060 18974 1116
rect 18974 1060 18978 1116
rect 18914 1056 18978 1060
rect 18994 1116 19058 1120
rect 18994 1060 18998 1116
rect 18998 1060 19054 1116
rect 19054 1060 19058 1116
rect 18994 1056 19058 1060
rect 24688 1116 24752 1120
rect 24688 1060 24692 1116
rect 24692 1060 24748 1116
rect 24748 1060 24752 1116
rect 24688 1056 24752 1060
rect 24768 1116 24832 1120
rect 24768 1060 24772 1116
rect 24772 1060 24828 1116
rect 24828 1060 24832 1116
rect 24768 1056 24832 1060
rect 24848 1116 24912 1120
rect 24848 1060 24852 1116
rect 24852 1060 24908 1116
rect 24908 1060 24912 1116
rect 24848 1056 24912 1060
rect 24928 1116 24992 1120
rect 24928 1060 24932 1116
rect 24932 1060 24988 1116
rect 24988 1060 24992 1116
rect 24928 1056 24992 1060
<< metal4 >>
rect 3911 8192 4231 8752
rect 3911 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4231 8192
rect 3911 7104 4231 8128
rect 3911 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4231 7104
rect 3911 6016 4231 7040
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 4928 4231 5952
rect 3911 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 2752 4231 3776
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3911 1664 4231 2688
rect 3911 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4231 1664
rect 3911 1040 4231 1600
rect 6878 8736 7198 8752
rect 6878 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7198 8736
rect 6878 7648 7198 8672
rect 6878 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7198 7648
rect 6878 6560 7198 7584
rect 6878 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7198 6560
rect 6878 5472 7198 6496
rect 6878 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7198 5472
rect 6878 4384 7198 5408
rect 6878 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7198 4384
rect 6878 3296 7198 4320
rect 6878 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7198 3296
rect 6878 2208 7198 3232
rect 6878 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7198 2208
rect 6878 1120 7198 2144
rect 6878 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7198 1120
rect 6878 1040 7198 1056
rect 9845 8192 10165 8752
rect 9845 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10165 8192
rect 9845 7104 10165 8128
rect 9845 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10165 7104
rect 9845 6016 10165 7040
rect 9845 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10165 6016
rect 9845 4928 10165 5952
rect 9845 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10165 4928
rect 9845 3840 10165 4864
rect 9845 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10165 3840
rect 9845 2752 10165 3776
rect 9845 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10165 2752
rect 9845 1664 10165 2688
rect 9845 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10165 1664
rect 9845 1040 10165 1600
rect 12812 8736 13132 8752
rect 12812 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13132 8736
rect 12812 7648 13132 8672
rect 12812 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13132 7648
rect 12812 6560 13132 7584
rect 12812 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13132 6560
rect 12812 5472 13132 6496
rect 12812 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13132 5472
rect 12812 4384 13132 5408
rect 12812 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13132 4384
rect 12812 3296 13132 4320
rect 12812 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13132 3296
rect 12812 2208 13132 3232
rect 12812 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13132 2208
rect 12812 1120 13132 2144
rect 12812 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13132 1120
rect 12812 1040 13132 1056
rect 15779 8192 16099 8752
rect 15779 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16099 8192
rect 15779 7104 16099 8128
rect 15779 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16099 7104
rect 15779 6016 16099 7040
rect 15779 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16099 6016
rect 15779 4928 16099 5952
rect 15779 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16099 4928
rect 15779 3840 16099 4864
rect 15779 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16099 3840
rect 15779 2752 16099 3776
rect 15779 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16099 2752
rect 15779 1664 16099 2688
rect 15779 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16099 1664
rect 15779 1040 16099 1600
rect 18746 8736 19066 8752
rect 18746 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19066 8736
rect 18746 7648 19066 8672
rect 18746 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19066 7648
rect 18746 6560 19066 7584
rect 18746 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19066 6560
rect 18746 5472 19066 6496
rect 18746 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19066 5472
rect 18746 4384 19066 5408
rect 18746 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19066 4384
rect 18746 3296 19066 4320
rect 18746 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19066 3296
rect 18746 2208 19066 3232
rect 18746 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19066 2208
rect 18746 1120 19066 2144
rect 18746 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19066 1120
rect 18746 1040 19066 1056
rect 21713 8192 22033 8752
rect 21713 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22033 8192
rect 21713 7104 22033 8128
rect 21713 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22033 7104
rect 21713 6016 22033 7040
rect 21713 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22033 6016
rect 21713 4928 22033 5952
rect 21713 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22033 4928
rect 21713 3840 22033 4864
rect 21713 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22033 3840
rect 21713 2752 22033 3776
rect 21713 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22033 2752
rect 21713 1664 22033 2688
rect 21713 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22033 1664
rect 21713 1040 22033 1600
rect 24680 8736 25000 8752
rect 24680 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 25000 8736
rect 24680 7648 25000 8672
rect 24680 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 25000 7648
rect 24680 6560 25000 7584
rect 24680 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25000 6560
rect 24680 5472 25000 6496
rect 24680 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25000 5472
rect 24680 4384 25000 5408
rect 24680 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25000 4384
rect 24680 3296 25000 4320
rect 24680 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25000 3296
rect 24680 2208 25000 3232
rect 24680 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25000 2208
rect 24680 1120 25000 2144
rect 24680 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 25000 1120
rect 24680 1040 25000 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3220 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_49
timestamp 1688980957
transform 1 0 5612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1688980957
transform 1 0 6072 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_72
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_78
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1688980957
transform 1 0 8648 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_88 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_148
timestamp 1688980957
transform 1 0 14720 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_152
timestamp 1688980957
transform 1 0 15088 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_161
timestamp 1688980957
transform 1 0 15916 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_175
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_184
timestamp 1688980957
transform 1 0 18032 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_188
timestamp 1688980957
transform 1 0 18400 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_200
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_206
timestamp 1688980957
transform 1 0 20056 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_210
timestamp 1688980957
transform 1 0 20424 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_218
timestamp 1688980957
transform 1 0 21160 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_231
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_239
timestamp 1688980957
transform 1 0 23092 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_75
timestamp 1688980957
transform 1 0 8004 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_83
timestamp 1688980957
transform 1 0 8740 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_88
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_96
timestamp 1688980957
transform 1 0 9936 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_100
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_104
timestamp 1688980957
transform 1 0 10672 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_116
timestamp 1688980957
transform 1 0 11776 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_124
timestamp 1688980957
transform 1 0 12512 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_131
timestamp 1688980957
transform 1 0 13156 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_135
timestamp 1688980957
transform 1 0 13524 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_142
timestamp 1688980957
transform 1 0 14168 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_153
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_158
timestamp 1688980957
transform 1 0 15640 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_162
timestamp 1688980957
transform 1 0 16008 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1688980957
transform 1 0 16376 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 1688980957
transform 1 0 18492 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_212
timestamp 1688980957
transform 1 0 20608 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_234
timestamp 1688980957
transform 1 0 22632 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_240
timestamp 1688980957
transform 1 0 23184 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_253
timestamp 1688980957
transform 1 0 24380 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_169
timestamp 1688980957
transform 1 0 16652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_173
timestamp 1688980957
transform 1 0 17020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_185
timestamp 1688980957
transform 1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_21
timestamp 1688980957
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_33
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_45
timestamp 1688980957
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_175
timestamp 1688980957
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_179
timestamp 1688980957
transform 1 0 17572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_191
timestamp 1688980957
transform 1 0 18676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_203
timestamp 1688980957
transform 1 0 19780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_215
timestamp 1688980957
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_241
timestamp 1688980957
transform 1 0 23276 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_254
timestamp 1688980957
transform 1 0 24472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_17
timestamp 1688980957
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1688980957
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_243
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_7
timestamp 1688980957
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_28
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_40
timestamp 1688980957
transform 1 0 4784 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_46
timestamp 1688980957
transform 1 0 5336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_63
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_67
timestamp 1688980957
transform 1 0 7268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_78
timestamp 1688980957
transform 1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_84
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_96
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_102
timestamp 1688980957
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_250
timestamp 1688980957
transform 1 0 24104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_254
timestamp 1688980957
transform 1 0 24472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_46
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_74
timestamp 1688980957
transform 1 0 7912 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_120
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_126
timestamp 1688980957
transform 1 0 12696 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_135
timestamp 1688980957
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_149
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_156
timestamp 1688980957
transform 1 0 15456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_184
timestamp 1688980957
transform 1 0 18032 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_207
timestamp 1688980957
transform 1 0 20148 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_243
timestamp 1688980957
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_7
timestamp 1688980957
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_26
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_36
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_64
timestamp 1688980957
transform 1 0 6992 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_94
timestamp 1688980957
transform 1 0 9752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_108
timestamp 1688980957
transform 1 0 11040 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_206
timestamp 1688980957
transform 1 0 20056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_247
timestamp 1688980957
transform 1 0 23828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_251
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 15364 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 16928 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 20148 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 21344 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 22540 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 23184 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 4600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 5796 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 10580 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 12420 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 13248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 14720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 14904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 19320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 19596 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 16100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 16376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 16652 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 16928 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  inst_clk_buf
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__00_
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__01_
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__02_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__03_
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__04_
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__05_
timestamp 1688980957
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__06_
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__07_
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__08_
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__09_
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__10_
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__11_
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__12_
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__13_
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__14_
timestamp 1688980957
transform 1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__15_
timestamp 1688980957
transform 1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__16_
timestamp 1688980957
transform 1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__17_
timestamp 1688980957
transform 1 0 9108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__18_
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__19_
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__20_
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__21_
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__22_
timestamp 1688980957
transform 1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__23_
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__24_
timestamp 1688980957
transform 1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__25_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__26_
timestamp 1688980957
transform 1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__27_
timestamp 1688980957
transform 1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__28_
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__29_
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__30_
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__31_
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__32_
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__33_
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__34_
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__35_
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform 1 0 21804 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 23368 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 23552 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output64
timestamp 1688980957
transform 1 0 23920 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output65
timestamp 1688980957
transform 1 0 23552 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output66
timestamp 1688980957
transform 1 0 23000 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 22448 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 21252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output70 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1688980957
transform 1 0 20884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 22172 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 22724 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output74
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 22356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 21896 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 22908 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 2944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 1840 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 1472 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 2392 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 1840 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 2024 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 2576 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1688980957
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 3956 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 4784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 5520 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1688980957
transform 1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 5888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1688980957
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 6440 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 6992 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 8096 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1688980957
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 24840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 14812 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 8372 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 12052 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 14444 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 15640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 16744 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 18124 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 20332 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 22816 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 23460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 15364 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 12880 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 10396 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 7728 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 10028 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 14904 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 16100 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 17296 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 18584 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 22356 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 23276 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 22080 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 23552 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 24104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 23828 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 14094 0 14150 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 15290 0 15346 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 17682 0 17738 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 18878 0 18934 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 21270 0 21326 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 22466 0 22522 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 24858 0 24914 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 3330 0 3386 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 4526 0 4582 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 6918 0 6974 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 8114 0 8170 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 10506 0 10562 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 11702 0 11758 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 20350 9840 20406 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 23110 9840 23166 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 23386 9840 23442 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 23662 9840 23718 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 23938 9840 23994 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 24214 9840 24270 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 24490 9840 24546 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 24766 9840 24822 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 25042 9840 25098 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 25318 9840 25374 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 25594 9840 25650 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 20626 9840 20682 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 20902 9840 20958 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 21178 9840 21234 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 21454 9840 21510 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 21730 9840 21786 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 22006 9840 22062 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 22282 9840 22338 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 22558 9840 22614 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 22834 9840 22890 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 202 9840 258 10000 0 FreeSans 224 90 0 0 N1BEG[0]
port 40 nsew signal tristate
flabel metal2 s 478 9840 534 10000 0 FreeSans 224 90 0 0 N1BEG[1]
port 41 nsew signal tristate
flabel metal2 s 754 9840 810 10000 0 FreeSans 224 90 0 0 N1BEG[2]
port 42 nsew signal tristate
flabel metal2 s 1030 9840 1086 10000 0 FreeSans 224 90 0 0 N1BEG[3]
port 43 nsew signal tristate
flabel metal2 s 1306 9840 1362 10000 0 FreeSans 224 90 0 0 N2BEG[0]
port 44 nsew signal tristate
flabel metal2 s 1582 9840 1638 10000 0 FreeSans 224 90 0 0 N2BEG[1]
port 45 nsew signal tristate
flabel metal2 s 1858 9840 1914 10000 0 FreeSans 224 90 0 0 N2BEG[2]
port 46 nsew signal tristate
flabel metal2 s 2134 9840 2190 10000 0 FreeSans 224 90 0 0 N2BEG[3]
port 47 nsew signal tristate
flabel metal2 s 2410 9840 2466 10000 0 FreeSans 224 90 0 0 N2BEG[4]
port 48 nsew signal tristate
flabel metal2 s 2686 9840 2742 10000 0 FreeSans 224 90 0 0 N2BEG[5]
port 49 nsew signal tristate
flabel metal2 s 2962 9840 3018 10000 0 FreeSans 224 90 0 0 N2BEG[6]
port 50 nsew signal tristate
flabel metal2 s 3238 9840 3294 10000 0 FreeSans 224 90 0 0 N2BEG[7]
port 51 nsew signal tristate
flabel metal2 s 3514 9840 3570 10000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 52 nsew signal tristate
flabel metal2 s 3790 9840 3846 10000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 53 nsew signal tristate
flabel metal2 s 4066 9840 4122 10000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 54 nsew signal tristate
flabel metal2 s 4342 9840 4398 10000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 55 nsew signal tristate
flabel metal2 s 4618 9840 4674 10000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 56 nsew signal tristate
flabel metal2 s 4894 9840 4950 10000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 57 nsew signal tristate
flabel metal2 s 5170 9840 5226 10000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 58 nsew signal tristate
flabel metal2 s 5446 9840 5502 10000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 59 nsew signal tristate
flabel metal2 s 5722 9840 5778 10000 0 FreeSans 224 90 0 0 N4BEG[0]
port 60 nsew signal tristate
flabel metal2 s 8482 9840 8538 10000 0 FreeSans 224 90 0 0 N4BEG[10]
port 61 nsew signal tristate
flabel metal2 s 8758 9840 8814 10000 0 FreeSans 224 90 0 0 N4BEG[11]
port 62 nsew signal tristate
flabel metal2 s 9034 9840 9090 10000 0 FreeSans 224 90 0 0 N4BEG[12]
port 63 nsew signal tristate
flabel metal2 s 9310 9840 9366 10000 0 FreeSans 224 90 0 0 N4BEG[13]
port 64 nsew signal tristate
flabel metal2 s 9586 9840 9642 10000 0 FreeSans 224 90 0 0 N4BEG[14]
port 65 nsew signal tristate
flabel metal2 s 9862 9840 9918 10000 0 FreeSans 224 90 0 0 N4BEG[15]
port 66 nsew signal tristate
flabel metal2 s 5998 9840 6054 10000 0 FreeSans 224 90 0 0 N4BEG[1]
port 67 nsew signal tristate
flabel metal2 s 6274 9840 6330 10000 0 FreeSans 224 90 0 0 N4BEG[2]
port 68 nsew signal tristate
flabel metal2 s 6550 9840 6606 10000 0 FreeSans 224 90 0 0 N4BEG[3]
port 69 nsew signal tristate
flabel metal2 s 6826 9840 6882 10000 0 FreeSans 224 90 0 0 N4BEG[4]
port 70 nsew signal tristate
flabel metal2 s 7102 9840 7158 10000 0 FreeSans 224 90 0 0 N4BEG[5]
port 71 nsew signal tristate
flabel metal2 s 7378 9840 7434 10000 0 FreeSans 224 90 0 0 N4BEG[6]
port 72 nsew signal tristate
flabel metal2 s 7654 9840 7710 10000 0 FreeSans 224 90 0 0 N4BEG[7]
port 73 nsew signal tristate
flabel metal2 s 7930 9840 7986 10000 0 FreeSans 224 90 0 0 N4BEG[8]
port 74 nsew signal tristate
flabel metal2 s 8206 9840 8262 10000 0 FreeSans 224 90 0 0 N4BEG[9]
port 75 nsew signal tristate
flabel metal2 s 10138 9840 10194 10000 0 FreeSans 224 90 0 0 S1END[0]
port 76 nsew signal input
flabel metal2 s 10414 9840 10470 10000 0 FreeSans 224 90 0 0 S1END[1]
port 77 nsew signal input
flabel metal2 s 10690 9840 10746 10000 0 FreeSans 224 90 0 0 S1END[2]
port 78 nsew signal input
flabel metal2 s 10966 9840 11022 10000 0 FreeSans 224 90 0 0 S1END[3]
port 79 nsew signal input
flabel metal2 s 11242 9840 11298 10000 0 FreeSans 224 90 0 0 S2END[0]
port 80 nsew signal input
flabel metal2 s 11518 9840 11574 10000 0 FreeSans 224 90 0 0 S2END[1]
port 81 nsew signal input
flabel metal2 s 11794 9840 11850 10000 0 FreeSans 224 90 0 0 S2END[2]
port 82 nsew signal input
flabel metal2 s 12070 9840 12126 10000 0 FreeSans 224 90 0 0 S2END[3]
port 83 nsew signal input
flabel metal2 s 12346 9840 12402 10000 0 FreeSans 224 90 0 0 S2END[4]
port 84 nsew signal input
flabel metal2 s 12622 9840 12678 10000 0 FreeSans 224 90 0 0 S2END[5]
port 85 nsew signal input
flabel metal2 s 12898 9840 12954 10000 0 FreeSans 224 90 0 0 S2END[6]
port 86 nsew signal input
flabel metal2 s 13174 9840 13230 10000 0 FreeSans 224 90 0 0 S2END[7]
port 87 nsew signal input
flabel metal2 s 13450 9840 13506 10000 0 FreeSans 224 90 0 0 S2MID[0]
port 88 nsew signal input
flabel metal2 s 13726 9840 13782 10000 0 FreeSans 224 90 0 0 S2MID[1]
port 89 nsew signal input
flabel metal2 s 14002 9840 14058 10000 0 FreeSans 224 90 0 0 S2MID[2]
port 90 nsew signal input
flabel metal2 s 14278 9840 14334 10000 0 FreeSans 224 90 0 0 S2MID[3]
port 91 nsew signal input
flabel metal2 s 14554 9840 14610 10000 0 FreeSans 224 90 0 0 S2MID[4]
port 92 nsew signal input
flabel metal2 s 14830 9840 14886 10000 0 FreeSans 224 90 0 0 S2MID[5]
port 93 nsew signal input
flabel metal2 s 15106 9840 15162 10000 0 FreeSans 224 90 0 0 S2MID[6]
port 94 nsew signal input
flabel metal2 s 15382 9840 15438 10000 0 FreeSans 224 90 0 0 S2MID[7]
port 95 nsew signal input
flabel metal2 s 15658 9840 15714 10000 0 FreeSans 224 90 0 0 S4END[0]
port 96 nsew signal input
flabel metal2 s 18418 9840 18474 10000 0 FreeSans 224 90 0 0 S4END[10]
port 97 nsew signal input
flabel metal2 s 18694 9840 18750 10000 0 FreeSans 224 90 0 0 S4END[11]
port 98 nsew signal input
flabel metal2 s 18970 9840 19026 10000 0 FreeSans 224 90 0 0 S4END[12]
port 99 nsew signal input
flabel metal2 s 19246 9840 19302 10000 0 FreeSans 224 90 0 0 S4END[13]
port 100 nsew signal input
flabel metal2 s 19522 9840 19578 10000 0 FreeSans 224 90 0 0 S4END[14]
port 101 nsew signal input
flabel metal2 s 19798 9840 19854 10000 0 FreeSans 224 90 0 0 S4END[15]
port 102 nsew signal input
flabel metal2 s 15934 9840 15990 10000 0 FreeSans 224 90 0 0 S4END[1]
port 103 nsew signal input
flabel metal2 s 16210 9840 16266 10000 0 FreeSans 224 90 0 0 S4END[2]
port 104 nsew signal input
flabel metal2 s 16486 9840 16542 10000 0 FreeSans 224 90 0 0 S4END[3]
port 105 nsew signal input
flabel metal2 s 16762 9840 16818 10000 0 FreeSans 224 90 0 0 S4END[4]
port 106 nsew signal input
flabel metal2 s 17038 9840 17094 10000 0 FreeSans 224 90 0 0 S4END[5]
port 107 nsew signal input
flabel metal2 s 17314 9840 17370 10000 0 FreeSans 224 90 0 0 S4END[6]
port 108 nsew signal input
flabel metal2 s 17590 9840 17646 10000 0 FreeSans 224 90 0 0 S4END[7]
port 109 nsew signal input
flabel metal2 s 17866 9840 17922 10000 0 FreeSans 224 90 0 0 S4END[8]
port 110 nsew signal input
flabel metal2 s 18142 9840 18198 10000 0 FreeSans 224 90 0 0 S4END[9]
port 111 nsew signal input
flabel metal2 s 938 0 994 160 0 FreeSans 224 90 0 0 UserCLK
port 112 nsew signal input
flabel metal2 s 20074 9840 20130 10000 0 FreeSans 224 90 0 0 UserCLKo
port 113 nsew signal tristate
flabel metal4 s 6878 1040 7198 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 12812 1040 13132 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 18746 1040 19066 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 24680 1040 25000 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 3911 1040 4231 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 9845 1040 10165 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 15779 1040 16099 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 21713 1040 22033 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
rlabel via1 13052 8704 13052 8704 0 VGND
rlabel metal1 12972 8160 12972 8160 0 VPWR
rlabel metal2 2215 68 2215 68 0 FrameStrobe[0]
rlabel metal2 14267 68 14267 68 0 FrameStrobe[10]
rlabel metal2 15463 68 15463 68 0 FrameStrobe[11]
rlabel metal2 16797 68 16797 68 0 FrameStrobe[12]
rlabel metal2 17855 68 17855 68 0 FrameStrobe[13]
rlabel metal2 19143 68 19143 68 0 FrameStrobe[14]
rlabel metal2 20247 68 20247 68 0 FrameStrobe[15]
rlabel metal2 21443 68 21443 68 0 FrameStrobe[16]
rlabel metal2 22639 68 22639 68 0 FrameStrobe[17]
rlabel metal2 23690 143 23690 143 0 FrameStrobe[18]
rlabel metal2 24886 398 24886 398 0 FrameStrobe[19]
rlabel metal2 3411 68 3411 68 0 FrameStrobe[1]
rlabel metal2 4699 68 4699 68 0 FrameStrobe[2]
rlabel metal2 5895 68 5895 68 0 FrameStrobe[3]
rlabel metal2 7229 68 7229 68 0 FrameStrobe[4]
rlabel metal2 8333 68 8333 68 0 FrameStrobe[5]
rlabel metal2 9529 68 9529 68 0 FrameStrobe[6]
rlabel metal2 10679 68 10679 68 0 FrameStrobe[7]
rlabel metal2 11875 68 11875 68 0 FrameStrobe[8]
rlabel metal2 12926 143 12926 143 0 FrameStrobe[9]
rlabel metal2 20378 9224 20378 9224 0 FrameStrobe_O[0]
rlabel metal2 23138 9224 23138 9224 0 FrameStrobe_O[10]
rlabel metal1 22816 7990 22816 7990 0 FrameStrobe_O[11]
rlabel metal2 23690 8952 23690 8952 0 FrameStrobe_O[12]
rlabel metal1 23874 6426 23874 6426 0 FrameStrobe_O[13]
rlabel metal1 24104 7514 24104 7514 0 FrameStrobe_O[14]
rlabel metal1 24426 6426 24426 6426 0 FrameStrobe_O[15]
rlabel metal1 24288 6834 24288 6834 0 FrameStrobe_O[16]
rlabel metal1 24242 7310 24242 7310 0 FrameStrobe_O[17]
rlabel metal1 24150 7446 24150 7446 0 FrameStrobe_O[18]
rlabel metal2 25622 8850 25622 8850 0 FrameStrobe_O[19]
rlabel metal2 20654 9224 20654 9224 0 FrameStrobe_O[1]
rlabel metal1 21528 8330 21528 8330 0 FrameStrobe_O[2]
rlabel metal1 21160 8058 21160 8058 0 FrameStrobe_O[3]
rlabel metal2 21482 9224 21482 9224 0 FrameStrobe_O[4]
rlabel metal2 21758 9462 21758 9462 0 FrameStrobe_O[5]
rlabel metal2 22034 9054 22034 9054 0 FrameStrobe_O[6]
rlabel metal2 22310 9309 22310 9309 0 FrameStrobe_O[7]
rlabel metal1 22448 7514 22448 7514 0 FrameStrobe_O[8]
rlabel metal2 22862 8952 22862 8952 0 FrameStrobe_O[9]
rlabel metal1 13708 1462 13708 1462 0 FrameStrobe_O_i\[0\]
rlabel metal1 14720 1530 14720 1530 0 FrameStrobe_O_i\[10\]
rlabel metal1 15916 1530 15916 1530 0 FrameStrobe_O_i\[11\]
rlabel metal1 17158 5882 17158 5882 0 FrameStrobe_O_i\[12\]
rlabel metal1 18400 1530 18400 1530 0 FrameStrobe_O_i\[13\]
rlabel metal1 22356 1462 22356 1462 0 FrameStrobe_O_i\[14\]
rlabel metal1 23506 1972 23506 1972 0 FrameStrobe_O_i\[15\]
rlabel metal2 22310 1734 22310 1734 0 FrameStrobe_O_i\[16\]
rlabel metal1 23230 1530 23230 1530 0 FrameStrobe_O_i\[17\]
rlabel metal1 24058 1530 24058 1530 0 FrameStrobe_O_i\[18\]
rlabel metal1 23782 1462 23782 1462 0 FrameStrobe_O_i\[19\]
rlabel metal1 14996 1190 14996 1190 0 FrameStrobe_O_i\[1\]
rlabel metal2 12926 1734 12926 1734 0 FrameStrobe_O_i\[2\]
rlabel metal1 10166 1530 10166 1530 0 FrameStrobe_O_i\[3\]
rlabel metal1 7498 1530 7498 1530 0 FrameStrobe_O_i\[4\]
rlabel metal1 8694 1530 8694 1530 0 FrameStrobe_O_i\[5\]
rlabel metal1 9706 1530 9706 1530 0 FrameStrobe_O_i\[6\]
rlabel metal1 11224 1530 11224 1530 0 FrameStrobe_O_i\[7\]
rlabel metal2 12650 1564 12650 1564 0 FrameStrobe_O_i\[8\]
rlabel metal1 13432 1530 13432 1530 0 FrameStrobe_O_i\[9\]
rlabel metal1 1288 6630 1288 6630 0 N1BEG[0]
rlabel metal2 506 9445 506 9445 0 N1BEG[1]
rlabel metal1 1196 6426 1196 6426 0 N1BEG[2]
rlabel metal1 1518 6834 1518 6834 0 N1BEG[3]
rlabel metal2 1334 8680 1334 8680 0 N2BEG[0]
rlabel metal2 1610 8952 1610 8952 0 N2BEG[1]
rlabel metal2 1886 9173 1886 9173 0 N2BEG[2]
rlabel metal2 2162 9445 2162 9445 0 N2BEG[3]
rlabel metal2 2438 8952 2438 8952 0 N2BEG[4]
rlabel metal2 2714 8952 2714 8952 0 N2BEG[5]
rlabel metal1 2898 8602 2898 8602 0 N2BEG[6]
rlabel metal2 3266 8952 3266 8952 0 N2BEG[7]
rlabel metal1 3358 7174 3358 7174 0 N2BEGb[0]
rlabel metal1 3680 7514 3680 7514 0 N2BEGb[1]
rlabel metal2 4094 9054 4094 9054 0 N2BEGb[2]
rlabel metal1 4324 8602 4324 8602 0 N2BEGb[3]
rlabel metal2 4646 8680 4646 8680 0 N2BEGb[4]
rlabel metal2 4922 8952 4922 8952 0 N2BEGb[5]
rlabel metal1 5014 8602 5014 8602 0 N2BEGb[6]
rlabel metal1 5428 8602 5428 8602 0 N2BEGb[7]
rlabel metal2 5750 9224 5750 9224 0 N4BEG[0]
rlabel metal1 8418 8602 8418 8602 0 N4BEG[10]
rlabel metal1 8740 8602 8740 8602 0 N4BEG[11]
rlabel metal1 9154 8602 9154 8602 0 N4BEG[12]
rlabel metal1 9476 8602 9476 8602 0 N4BEG[13]
rlabel metal2 9614 9088 9614 9088 0 N4BEG[14]
rlabel metal1 10902 8364 10902 8364 0 N4BEG[15]
rlabel metal2 6026 8952 6026 8952 0 N4BEG[1]
rlabel metal1 6026 7990 6026 7990 0 N4BEG[2]
rlabel metal2 6578 8952 6578 8952 0 N4BEG[3]
rlabel metal1 6716 8602 6716 8602 0 N4BEG[4]
rlabel metal2 7130 9326 7130 9326 0 N4BEG[5]
rlabel metal1 7590 8058 7590 8058 0 N4BEG[6]
rlabel metal1 7544 8602 7544 8602 0 N4BEG[7]
rlabel metal1 7958 8602 7958 8602 0 N4BEG[8]
rlabel metal2 8234 9190 8234 9190 0 N4BEG[9]
rlabel metal2 10166 9241 10166 9241 0 S1END[0]
rlabel metal2 10442 8850 10442 8850 0 S1END[1]
rlabel metal2 10718 8850 10718 8850 0 S1END[2]
rlabel metal2 10994 8850 10994 8850 0 S1END[3]
rlabel metal2 11270 9173 11270 9173 0 S2END[0]
rlabel metal2 11546 9377 11546 9377 0 S2END[1]
rlabel metal2 11822 9377 11822 9377 0 S2END[2]
rlabel metal2 12098 9156 12098 9156 0 S2END[3]
rlabel metal2 12374 9377 12374 9377 0 S2END[4]
rlabel metal2 12650 9564 12650 9564 0 S2END[5]
rlabel metal2 12926 9377 12926 9377 0 S2END[6]
rlabel metal2 13202 9445 13202 9445 0 S2END[7]
rlabel metal2 13478 9156 13478 9156 0 S2MID[0]
rlabel metal2 13754 9156 13754 9156 0 S2MID[1]
rlabel metal2 14030 9190 14030 9190 0 S2MID[2]
rlabel metal2 14306 9836 14306 9836 0 S2MID[3]
rlabel metal2 14582 9122 14582 9122 0 S2MID[4]
rlabel metal2 14858 8850 14858 8850 0 S2MID[5]
rlabel metal2 15134 8850 15134 8850 0 S2MID[6]
rlabel metal2 15410 9088 15410 9088 0 S2MID[7]
rlabel metal2 15686 9377 15686 9377 0 S4END[0]
rlabel metal2 18446 9105 18446 9105 0 S4END[10]
rlabel metal2 18722 9496 18722 9496 0 S4END[11]
rlabel metal2 18998 9513 18998 9513 0 S4END[12]
rlabel metal2 19274 8850 19274 8850 0 S4END[13]
rlabel metal2 19550 8850 19550 8850 0 S4END[14]
rlabel metal2 19826 8850 19826 8850 0 S4END[15]
rlabel metal2 15962 9377 15962 9377 0 S4END[1]
rlabel metal2 16238 8884 16238 8884 0 S4END[2]
rlabel metal2 16514 8918 16514 8918 0 S4END[3]
rlabel metal2 16790 8816 16790 8816 0 S4END[4]
rlabel metal2 17066 8884 17066 8884 0 S4END[5]
rlabel metal2 17342 8918 17342 8918 0 S4END[6]
rlabel metal2 17618 9224 17618 9224 0 S4END[7]
rlabel metal2 17894 9173 17894 9173 0 S4END[8]
rlabel metal2 18170 8850 18170 8850 0 S4END[9]
rlabel metal2 966 704 966 704 0 UserCLK
rlabel metal1 20240 8602 20240 8602 0 UserCLKo
rlabel metal1 2438 748 2438 748 0 net1
rlabel metal1 24012 1326 24012 1326 0 net10
rlabel metal2 17250 8772 17250 8772 0 net100
rlabel metal2 16974 8806 16974 8806 0 net101
rlabel metal2 16698 8840 16698 8840 0 net102
rlabel metal1 14858 7990 14858 7990 0 net103
rlabel metal2 15870 8738 15870 8738 0 net104
rlabel metal2 5474 7650 5474 7650 0 net105
rlabel metal1 5934 7514 5934 7514 0 net106
rlabel metal1 6624 7514 6624 7514 0 net107
rlabel metal1 18906 7990 18906 7990 0 net108
rlabel metal2 18078 7344 18078 7344 0 net109
rlabel metal1 23690 1292 23690 1292 0 net11
rlabel metal1 18860 8602 18860 8602 0 net110
rlabel metal1 17940 8058 17940 8058 0 net111
rlabel metal2 18262 8976 18262 8976 0 net112
rlabel metal1 17204 8330 17204 8330 0 net113
rlabel metal2 16882 1088 16882 1088 0 net114
rlabel metal1 3634 1224 3634 1224 0 net12
rlabel metal2 4646 1088 4646 1088 0 net13
rlabel metal2 5842 1020 5842 1020 0 net14
rlabel metal1 7452 1326 7452 1326 0 net15
rlabel metal1 8786 1326 8786 1326 0 net16
rlabel metal1 9798 1292 9798 1292 0 net17
rlabel metal1 11086 1292 11086 1292 0 net18
rlabel metal1 12282 1292 12282 1292 0 net19
rlabel metal1 14674 1292 14674 1292 0 net2
rlabel metal1 13386 1292 13386 1292 0 net20
rlabel metal1 9982 7514 9982 7514 0 net21
rlabel metal1 6578 7344 6578 7344 0 net22
rlabel metal1 7682 7310 7682 7310 0 net23
rlabel metal1 7958 7344 7958 7344 0 net24
rlabel metal1 8464 7378 8464 7378 0 net25
rlabel metal1 9568 7378 9568 7378 0 net26
rlabel metal1 9338 7820 9338 7820 0 net27
rlabel metal2 9706 8245 9706 8245 0 net28
rlabel metal1 12282 7888 12282 7888 0 net29
rlabel metal1 15870 1292 15870 1292 0 net3
rlabel metal1 11362 7854 11362 7854 0 net30
rlabel metal2 13018 8211 13018 8211 0 net31
rlabel metal1 12926 7990 12926 7990 0 net32
rlabel metal1 11730 8398 11730 8398 0 net33
rlabel metal1 12282 8432 12282 8432 0 net34
rlabel metal1 12650 8500 12650 8500 0 net35
rlabel metal1 12834 8466 12834 8466 0 net36
rlabel metal1 13754 8398 13754 8398 0 net37
rlabel metal1 14582 8058 14582 8058 0 net38
rlabel metal2 15226 8262 15226 8262 0 net39
rlabel metal1 16974 1258 16974 1258 0 net4
rlabel metal1 15594 8500 15594 8500 0 net40
rlabel metal1 15778 8058 15778 8058 0 net41
rlabel metal1 18538 7820 18538 7820 0 net42
rlabel metal1 18814 7888 18814 7888 0 net43
rlabel metal2 20010 9078 20010 9078 0 net44
rlabel metal2 19550 7497 19550 7497 0 net45
rlabel metal2 19826 7582 19826 7582 0 net46
rlabel metal2 20102 7565 20102 7565 0 net47
rlabel metal1 15778 7888 15778 7888 0 net48
rlabel metal1 16652 8058 16652 8058 0 net49
rlabel metal1 18354 1292 18354 1292 0 net5
rlabel metal2 16698 8058 16698 8058 0 net50
rlabel metal1 17204 8058 17204 8058 0 net51
rlabel metal2 17250 8194 17250 8194 0 net52
rlabel metal1 17664 8058 17664 8058 0 net53
rlabel metal1 18216 8466 18216 8466 0 net54
rlabel metal1 17940 7854 17940 7854 0 net55
rlabel metal1 18492 7990 18492 7990 0 net56
rlabel metal1 1610 952 1610 952 0 net57
rlabel metal1 15226 1802 15226 1802 0 net58
rlabel metal1 22954 2584 22954 2584 0 net59
rlabel metal1 22218 1326 22218 1326 0 net6
rlabel metal1 17066 2074 17066 2074 0 net60
rlabel metal2 23874 6936 23874 6936 0 net61
rlabel metal1 23506 1836 23506 1836 0 net62
rlabel metal2 22402 2244 22402 2244 0 net63
rlabel metal1 23368 1734 23368 1734 0 net64
rlabel metal2 22126 4420 22126 4420 0 net65
rlabel metal1 23368 2074 23368 2074 0 net66
rlabel metal2 24150 2210 24150 2210 0 net67
rlabel metal1 23828 2074 23828 2074 0 net68
rlabel metal1 18216 1734 18216 1734 0 net69
rlabel metal1 20378 1530 20378 1530 0 net7
rlabel metal1 13432 2074 13432 2074 0 net70
rlabel metal2 10626 2176 10626 2176 0 net71
rlabel metal2 22264 7684 22264 7684 0 net72
rlabel metal2 22310 4572 22310 4572 0 net73
rlabel metal2 23046 4539 23046 4539 0 net74
rlabel metal2 22494 5151 22494 5151 0 net75
rlabel metal1 12834 2040 12834 2040 0 net76
rlabel metal1 22862 7786 22862 7786 0 net77
rlabel metal2 7774 7106 7774 7106 0 net78
rlabel metal2 7498 7922 7498 7922 0 net79
rlabel metal1 21850 1326 21850 1326 0 net8
rlabel metal2 6394 6766 6394 6766 0 net80
rlabel metal2 9798 7310 9798 7310 0 net81
rlabel metal2 1978 7633 1978 7633 0 net82
rlabel metal2 1794 8500 1794 8500 0 net83
rlabel metal2 2714 7701 2714 7701 0 net84
rlabel metal1 1978 8432 1978 8432 0 net85
rlabel metal2 2346 8534 2346 8534 0 net86
rlabel metal1 13202 8262 13202 8262 0 net87
rlabel metal1 11776 8602 11776 8602 0 net88
rlabel metal1 3266 7786 3266 7786 0 net89
rlabel metal1 23046 1292 23046 1292 0 net9
rlabel metal1 2990 7344 2990 7344 0 net90
rlabel metal1 3864 7378 3864 7378 0 net91
rlabel metal1 4692 7854 4692 7854 0 net92
rlabel metal1 9614 7718 9614 7718 0 net93
rlabel metal1 4922 7378 4922 7378 0 net94
rlabel metal1 4922 7752 4922 7752 0 net95
rlabel metal1 8648 7514 8648 7514 0 net96
rlabel metal1 7958 7514 7958 7514 0 net97
rlabel metal1 5704 7514 5704 7514 0 net98
rlabel metal2 17526 8908 17526 8908 0 net99
<< properties >>
string FIXED_BBOX 0 0 26000 10000
<< end >>
