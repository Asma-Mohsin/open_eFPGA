magic
tech sky130A
magscale 1 2
timestamp 1733308638
<< viali >>
rect 1593 43401 1627 43435
rect 2329 43401 2363 43435
rect 2881 43401 2915 43435
rect 3433 43401 3467 43435
rect 3985 43401 4019 43435
rect 4537 43401 4571 43435
rect 5273 43401 5307 43435
rect 5917 43401 5951 43435
rect 6745 43401 6779 43435
rect 7481 43401 7515 43435
rect 8217 43401 8251 43435
rect 9137 43401 9171 43435
rect 9689 43401 9723 43435
rect 10425 43401 10459 43435
rect 11713 43401 11747 43435
rect 12265 43401 12299 43435
rect 12633 43401 12667 43435
rect 13277 43401 13311 43435
rect 13829 43401 13863 43435
rect 1501 43265 1535 43299
rect 2145 43265 2179 43299
rect 2789 43265 2823 43299
rect 3249 43265 3283 43299
rect 3801 43265 3835 43299
rect 4445 43265 4479 43299
rect 5089 43265 5123 43299
rect 5825 43265 5859 43299
rect 6653 43265 6687 43299
rect 7297 43265 7331 43299
rect 8125 43265 8159 43299
rect 8953 43265 8987 43299
rect 9597 43265 9631 43299
rect 10241 43265 10275 43299
rect 11621 43265 11655 43299
rect 12081 43265 12115 43299
rect 12541 43265 12575 43299
rect 13093 43265 13127 43299
rect 13553 43265 13587 43299
rect 14289 43265 14323 43299
rect 14105 43061 14139 43095
rect 2881 42857 2915 42891
rect 3341 42857 3375 42891
rect 4169 42857 4203 42891
rect 4905 42857 4939 42891
rect 5641 42857 5675 42891
rect 6377 42857 6411 42891
rect 7113 42857 7147 42891
rect 7849 42857 7883 42891
rect 8585 42857 8619 42891
rect 9229 42857 9263 42891
rect 10241 42857 10275 42891
rect 10793 42857 10827 42891
rect 12265 42857 12299 42891
rect 13001 42857 13035 42891
rect 11529 42789 11563 42823
rect 13829 42721 13863 42755
rect 3525 42653 3559 42687
rect 4353 42653 4387 42687
rect 5089 42653 5123 42687
rect 5825 42653 5859 42687
rect 6561 42653 6595 42687
rect 7297 42653 7331 42687
rect 8033 42653 8067 42687
rect 8769 42653 8803 42687
rect 9413 42653 9447 42687
rect 10057 42653 10091 42687
rect 10977 42653 11011 42687
rect 11713 42653 11747 42687
rect 12449 42653 12483 42687
rect 13185 42653 13219 42687
rect 14289 42653 14323 42687
rect 1409 42585 1443 42619
rect 13553 42585 13587 42619
rect 9689 42517 9723 42551
rect 14105 42517 14139 42551
rect 2053 42313 2087 42347
rect 4077 42313 4111 42347
rect 4905 42313 4939 42347
rect 13737 42313 13771 42347
rect 14197 42313 14231 42347
rect 14105 42245 14139 42279
rect 2237 42177 2271 42211
rect 4261 42177 4295 42211
rect 5089 42177 5123 42211
rect 13921 42177 13955 42211
rect 1409 41089 1443 41123
rect 1593 40885 1627 40919
rect 1409 40477 1443 40511
rect 13553 40409 13587 40443
rect 1593 40341 1627 40375
rect 13829 40341 13863 40375
rect 9229 40137 9263 40171
rect 10057 40137 10091 40171
rect 9413 40001 9447 40035
rect 10241 40001 10275 40035
rect 13369 40001 13403 40035
rect 13921 40001 13955 40035
rect 13645 39797 13679 39831
rect 14197 39797 14231 39831
rect 13001 39593 13035 39627
rect 8953 39525 8987 39559
rect 9505 39525 9539 39559
rect 1409 39389 1443 39423
rect 9137 39389 9171 39423
rect 9689 39389 9723 39423
rect 12909 39389 12943 39423
rect 13185 39389 13219 39423
rect 14197 39389 14231 39423
rect 13553 39321 13587 39355
rect 13921 39321 13955 39355
rect 1593 39253 1627 39287
rect 12725 39253 12759 39287
rect 14381 39253 14415 39287
rect 12725 39049 12759 39083
rect 1409 38913 1443 38947
rect 12909 38913 12943 38947
rect 13185 38913 13219 38947
rect 13369 38913 13403 38947
rect 13921 38913 13955 38947
rect 13001 38777 13035 38811
rect 1593 38709 1627 38743
rect 13645 38709 13679 38743
rect 14197 38709 14231 38743
rect 12725 38505 12759 38539
rect 12449 38437 12483 38471
rect 12633 38301 12667 38335
rect 12909 38301 12943 38335
rect 13185 38301 13219 38335
rect 13461 38301 13495 38335
rect 13645 38301 13679 38335
rect 14197 38301 14231 38335
rect 13001 38165 13035 38199
rect 13277 38165 13311 38199
rect 13829 38165 13863 38199
rect 14381 38165 14415 38199
rect 11529 37961 11563 37995
rect 11805 37961 11839 37995
rect 1409 37825 1443 37859
rect 11713 37825 11747 37859
rect 11989 37825 12023 37859
rect 12817 37825 12851 37859
rect 13001 37825 13035 37859
rect 13369 37825 13403 37859
rect 13553 37825 13587 37859
rect 14105 37825 14139 37859
rect 1593 37689 1627 37723
rect 12633 37621 12667 37655
rect 13829 37621 13863 37655
rect 14381 37621 14415 37655
rect 10793 37417 10827 37451
rect 12633 37417 12667 37451
rect 13185 37417 13219 37451
rect 12909 37349 12943 37383
rect 1777 37281 1811 37315
rect 13829 37281 13863 37315
rect 10977 37213 11011 37247
rect 12541 37213 12575 37247
rect 12817 37213 12851 37247
rect 13093 37213 13127 37247
rect 13369 37213 13403 37247
rect 14197 37213 14231 37247
rect 1501 37145 1535 37179
rect 13553 37145 13587 37179
rect 12357 37077 12391 37111
rect 14381 37077 14415 37111
rect 11897 36873 11931 36907
rect 12725 36873 12759 36907
rect 14381 36873 14415 36907
rect 12081 36737 12115 36771
rect 12357 36737 12391 36771
rect 12633 36737 12667 36771
rect 12909 36737 12943 36771
rect 13185 36737 13219 36771
rect 13553 36737 13587 36771
rect 13921 36737 13955 36771
rect 14105 36737 14139 36771
rect 12173 36601 12207 36635
rect 12449 36533 12483 36567
rect 13737 36533 13771 36567
rect 9137 36329 9171 36363
rect 11529 36329 11563 36363
rect 12357 36329 12391 36363
rect 12633 36329 12667 36363
rect 11805 36261 11839 36295
rect 9321 36125 9355 36159
rect 11713 36125 11747 36159
rect 11989 36125 12023 36159
rect 12265 36125 12299 36159
rect 12541 36125 12575 36159
rect 12817 36125 12851 36159
rect 14197 36125 14231 36159
rect 1501 36057 1535 36091
rect 1869 36057 1903 36091
rect 13001 36057 13035 36091
rect 13553 36057 13587 36091
rect 13921 36057 13955 36091
rect 12081 35989 12115 36023
rect 13277 35989 13311 36023
rect 14381 35989 14415 36023
rect 1777 35785 1811 35819
rect 8401 35785 8435 35819
rect 10149 35785 10183 35819
rect 11529 35785 11563 35819
rect 11805 35785 11839 35819
rect 12449 35717 12483 35751
rect 13001 35717 13035 35751
rect 1409 35649 1443 35683
rect 1961 35649 1995 35683
rect 8585 35649 8619 35683
rect 10333 35649 10367 35683
rect 11345 35649 11379 35683
rect 11713 35649 11747 35683
rect 11989 35649 12023 35683
rect 12265 35649 12299 35683
rect 13369 35649 13403 35683
rect 13553 35649 13587 35683
rect 14105 35649 14139 35683
rect 11161 35513 11195 35547
rect 12081 35513 12115 35547
rect 1593 35445 1627 35479
rect 12725 35445 12759 35479
rect 13829 35445 13863 35479
rect 14381 35445 14415 35479
rect 1593 35241 1627 35275
rect 9321 35241 9355 35275
rect 11253 35241 11287 35275
rect 14105 35173 14139 35207
rect 11529 35105 11563 35139
rect 1777 35037 1811 35071
rect 9505 35037 9539 35071
rect 11437 35037 11471 35071
rect 11771 35037 11805 35071
rect 13001 35037 13035 35071
rect 14289 35037 14323 35071
rect 13553 34969 13587 35003
rect 13921 34969 13955 35003
rect 12541 34901 12575 34935
rect 13277 34901 13311 34935
rect 1593 34697 1627 34731
rect 10425 34697 10459 34731
rect 10701 34697 10735 34731
rect 10977 34697 11011 34731
rect 11529 34697 11563 34731
rect 11897 34629 11931 34663
rect 13001 34629 13035 34663
rect 1409 34561 1443 34595
rect 10609 34561 10643 34595
rect 10885 34561 10919 34595
rect 11161 34561 11195 34595
rect 11713 34561 11747 34595
rect 12265 34561 12299 34595
rect 12449 34561 12483 34595
rect 13369 34561 13403 34595
rect 13553 34561 13587 34595
rect 14105 34561 14139 34595
rect 14473 34561 14507 34595
rect 12725 34493 12759 34527
rect 13829 34357 13863 34391
rect 10241 34153 10275 34187
rect 10517 34153 10551 34187
rect 12173 34017 12207 34051
rect 1409 33949 1443 33983
rect 10425 33949 10459 33983
rect 10701 33949 10735 33983
rect 10793 33949 10827 33983
rect 11067 33949 11101 33983
rect 12415 33939 12449 33973
rect 13737 33949 13771 33983
rect 14289 33949 14323 33983
rect 1593 33813 1627 33847
rect 11805 33813 11839 33847
rect 13185 33813 13219 33847
rect 13553 33813 13587 33847
rect 14105 33813 14139 33847
rect 11621 33609 11655 33643
rect 13553 33541 13587 33575
rect 11805 33473 11839 33507
rect 12171 33473 12205 33507
rect 14105 33473 14139 33507
rect 11897 33405 11931 33439
rect 12909 33269 12943 33303
rect 13829 33269 13863 33303
rect 14197 33269 14231 33303
rect 9505 33065 9539 33099
rect 10517 33065 10551 33099
rect 11253 33065 11287 33099
rect 14105 33065 14139 33099
rect 9965 32997 9999 33031
rect 10977 32997 11011 33031
rect 12725 32929 12759 32963
rect 1409 32861 1443 32895
rect 9689 32861 9723 32895
rect 10149 32861 10183 32895
rect 10701 32861 10735 32895
rect 11161 32861 11195 32895
rect 11437 32861 11471 32895
rect 11713 32861 11747 32895
rect 13001 32861 13035 32895
rect 14289 32861 14323 32895
rect 11897 32793 11931 32827
rect 12449 32793 12483 32827
rect 13369 32793 13403 32827
rect 13553 32793 13587 32827
rect 13921 32793 13955 32827
rect 1593 32725 1627 32759
rect 11529 32725 11563 32759
rect 12173 32725 12207 32759
rect 2053 32521 2087 32555
rect 1409 32385 1443 32419
rect 2237 32385 2271 32419
rect 7021 32385 7055 32419
rect 7279 32415 7313 32449
rect 8401 32385 8435 32419
rect 8659 32415 8693 32449
rect 10299 32385 10333 32419
rect 11771 32385 11805 32419
rect 13001 32385 13035 32419
rect 13553 32385 13587 32419
rect 13921 32385 13955 32419
rect 14105 32385 14139 32419
rect 10057 32317 10091 32351
rect 11529 32317 11563 32351
rect 11069 32249 11103 32283
rect 1593 32181 1627 32215
rect 8033 32181 8067 32215
rect 9413 32181 9447 32215
rect 12541 32181 12575 32215
rect 13277 32181 13311 32215
rect 14381 32181 14415 32215
rect 8953 31977 8987 32011
rect 10517 31977 10551 32011
rect 10793 31977 10827 32011
rect 11069 31977 11103 32011
rect 14105 31977 14139 32011
rect 12639 31841 12673 31875
rect 13829 31841 13863 31875
rect 9137 31773 9171 31807
rect 10701 31773 10735 31807
rect 10977 31773 11011 31807
rect 11253 31773 11287 31807
rect 11529 31773 11563 31807
rect 11897 31773 11931 31807
rect 11989 31773 12023 31807
rect 12173 31773 12207 31807
rect 12909 31773 12943 31807
rect 13047 31773 13081 31807
rect 13185 31773 13219 31807
rect 14289 31773 14323 31807
rect 10701 31433 10735 31467
rect 10977 31433 11011 31467
rect 13369 31365 13403 31399
rect 13553 31365 13587 31399
rect 1409 31297 1443 31331
rect 9321 31297 9355 31331
rect 9595 31297 9629 31331
rect 10885 31297 10919 31331
rect 11161 31297 11195 31331
rect 11713 31297 11747 31331
rect 12725 31297 12759 31331
rect 14105 31297 14139 31331
rect 11529 31229 11563 31263
rect 12173 31229 12207 31263
rect 12449 31229 12483 31263
rect 12566 31229 12600 31263
rect 1593 31093 1627 31127
rect 10333 31093 10367 31127
rect 13829 31093 13863 31127
rect 14381 31093 14415 31127
rect 13921 30889 13955 30923
rect 12725 30821 12759 30855
rect 7205 30753 7239 30787
rect 11345 30753 11379 30787
rect 13001 30753 13035 30787
rect 13277 30753 13311 30787
rect 1409 30685 1443 30719
rect 7463 30655 7497 30689
rect 11621 30685 11655 30719
rect 12081 30685 12115 30719
rect 12265 30685 12299 30719
rect 13139 30685 13173 30719
rect 11069 30617 11103 30651
rect 11989 30617 12023 30651
rect 1593 30549 1627 30583
rect 8217 30549 8251 30583
rect 10057 30277 10091 30311
rect 10977 30277 11011 30311
rect 11345 30277 11379 30311
rect 6837 30209 6871 30243
rect 7111 30209 7145 30243
rect 9413 30209 9447 30243
rect 10425 30209 10459 30243
rect 11805 30209 11839 30243
rect 12171 30209 12205 30243
rect 13553 30209 13587 30243
rect 13921 30209 13955 30243
rect 14105 30209 14139 30243
rect 8217 30141 8251 30175
rect 8401 30141 8435 30175
rect 9137 30141 9171 30175
rect 9275 30141 9309 30175
rect 11897 30141 11931 30175
rect 7849 30073 7883 30107
rect 8861 30073 8895 30107
rect 11621 30073 11655 30107
rect 10701 30005 10735 30039
rect 12909 30005 12943 30039
rect 14381 30005 14415 30039
rect 12725 29801 12759 29835
rect 11345 29733 11379 29767
rect 8953 29665 8987 29699
rect 1409 29597 1443 29631
rect 9227 29587 9261 29621
rect 10333 29597 10367 29631
rect 10607 29597 10641 29631
rect 11713 29597 11747 29631
rect 11987 29597 12021 29631
rect 13553 29529 13587 29563
rect 1593 29461 1627 29495
rect 9965 29461 9999 29495
rect 13645 29461 13679 29495
rect 9873 29257 9907 29291
rect 11529 29189 11563 29223
rect 13921 29189 13955 29223
rect 1409 29121 1443 29155
rect 8217 29121 8251 29155
rect 9229 29121 9263 29155
rect 10331 29131 10365 29165
rect 12173 29121 12207 29155
rect 13737 29121 13771 29155
rect 8033 29053 8067 29087
rect 8677 29053 8711 29087
rect 8953 29053 8987 29087
rect 9091 29053 9125 29087
rect 10057 29053 10091 29087
rect 12311 29053 12345 29087
rect 12449 29053 12483 29087
rect 12725 29053 12759 29087
rect 13185 29053 13219 29087
rect 13369 29053 13403 29087
rect 1593 28985 1627 29019
rect 14197 28985 14231 29019
rect 11069 28917 11103 28951
rect 11069 28713 11103 28747
rect 13921 28713 13955 28747
rect 9873 28645 9907 28679
rect 12725 28645 12759 28679
rect 6377 28577 6411 28611
rect 9413 28577 9447 28611
rect 10149 28577 10183 28611
rect 10425 28577 10459 28611
rect 12265 28577 12299 28611
rect 13139 28577 13173 28611
rect 13277 28577 13311 28611
rect 6651 28509 6685 28543
rect 9229 28509 9263 28543
rect 10287 28509 10321 28543
rect 12081 28509 12115 28543
rect 13001 28509 13035 28543
rect 11621 28441 11655 28475
rect 7389 28373 7423 28407
rect 11897 28373 11931 28407
rect 1593 28169 1627 28203
rect 10517 28169 10551 28203
rect 1409 28033 1443 28067
rect 7297 28033 7331 28067
rect 7555 28063 7589 28097
rect 8677 28033 8711 28067
rect 9735 28033 9769 28067
rect 12063 28043 12097 28077
rect 13185 28033 13219 28067
rect 13427 28033 13461 28067
rect 8861 27965 8895 27999
rect 9597 27965 9631 27999
rect 9873 27965 9907 27999
rect 11805 27965 11839 27999
rect 8309 27897 8343 27931
rect 9321 27897 9355 27931
rect 12817 27829 12851 27863
rect 14197 27829 14231 27863
rect 9965 27625 9999 27659
rect 5917 27557 5951 27591
rect 6929 27557 6963 27591
rect 6469 27489 6503 27523
rect 7205 27489 7239 27523
rect 7322 27489 7356 27523
rect 8953 27489 8987 27523
rect 12633 27489 12667 27523
rect 4905 27421 4939 27455
rect 5163 27391 5197 27425
rect 6285 27421 6319 27455
rect 7481 27421 7515 27455
rect 9195 27421 9229 27455
rect 11989 27421 12023 27455
rect 12907 27421 12941 27455
rect 1501 27353 1535 27387
rect 8125 27353 8159 27387
rect 10885 27353 10919 27387
rect 11437 27353 11471 27387
rect 12357 27353 12391 27387
rect 1593 27285 1627 27319
rect 11161 27285 11195 27319
rect 11713 27285 11747 27319
rect 13645 27285 13679 27319
rect 2973 27081 3007 27115
rect 8585 27081 8619 27115
rect 13369 27013 13403 27047
rect 13737 27013 13771 27047
rect 2789 26945 2823 26979
rect 5147 26945 5181 26979
rect 10207 26945 10241 26979
rect 11529 26945 11563 26979
rect 12449 26945 12483 26979
rect 12725 26945 12759 26979
rect 4905 26877 4939 26911
rect 6745 26877 6779 26911
rect 6929 26877 6963 26911
rect 7665 26877 7699 26911
rect 7782 26877 7816 26911
rect 7941 26877 7975 26911
rect 9965 26877 9999 26911
rect 11713 26877 11747 26911
rect 12587 26877 12621 26911
rect 5917 26809 5951 26843
rect 7389 26809 7423 26843
rect 10977 26809 11011 26843
rect 12173 26809 12207 26843
rect 14013 26741 14047 26775
rect 2881 26537 2915 26571
rect 7757 26537 7791 26571
rect 11529 26537 11563 26571
rect 13921 26537 13955 26571
rect 1685 26469 1719 26503
rect 12725 26469 12759 26503
rect 6745 26401 6779 26435
rect 13001 26401 13035 26435
rect 13277 26401 13311 26435
rect 3065 26333 3099 26367
rect 6987 26333 7021 26367
rect 10517 26333 10551 26367
rect 10759 26333 10793 26367
rect 12081 26333 12115 26367
rect 12265 26333 12299 26367
rect 13139 26333 13173 26367
rect 1501 26265 1535 26299
rect 14473 25993 14507 26027
rect 12173 25925 12207 25959
rect 1685 25857 1719 25891
rect 9871 25857 9905 25891
rect 11621 25857 11655 25891
rect 12817 25857 12851 25891
rect 13691 25857 13725 25891
rect 13829 25857 13863 25891
rect 1409 25789 1443 25823
rect 9597 25789 9631 25823
rect 12633 25789 12667 25823
rect 13553 25789 13587 25823
rect 13277 25721 13311 25755
rect 10609 25653 10643 25687
rect 11897 25653 11931 25687
rect 12449 25653 12483 25687
rect 10793 25449 10827 25483
rect 13001 25449 13035 25483
rect 8493 25381 8527 25415
rect 9597 25381 9631 25415
rect 10149 25313 10183 25347
rect 11989 25313 12023 25347
rect 7481 25245 7515 25279
rect 7755 25245 7789 25279
rect 8953 25245 8987 25279
rect 9137 25245 9171 25279
rect 9873 25245 9907 25279
rect 9990 25245 10024 25279
rect 12231 25245 12265 25279
rect 11529 25177 11563 25211
rect 11897 25177 11931 25211
rect 13553 25177 13587 25211
rect 13921 25177 13955 25211
rect 9505 24905 9539 24939
rect 1501 24769 1535 24803
rect 6743 24769 6777 24803
rect 8735 24769 8769 24803
rect 10331 24769 10365 24803
rect 11771 24769 11805 24803
rect 13183 24769 13217 24803
rect 6469 24701 6503 24735
rect 8493 24701 8527 24735
rect 10057 24701 10091 24735
rect 11529 24701 11563 24735
rect 12909 24701 12943 24735
rect 1685 24633 1719 24667
rect 7481 24565 7515 24599
rect 11069 24565 11103 24599
rect 12541 24565 12575 24599
rect 13921 24565 13955 24599
rect 9965 24361 9999 24395
rect 12633 24361 12667 24395
rect 7573 24293 7607 24327
rect 11437 24293 11471 24327
rect 7966 24225 8000 24259
rect 8125 24225 8159 24259
rect 11713 24225 11747 24259
rect 11851 24225 11885 24259
rect 11989 24225 12023 24259
rect 5549 24157 5583 24191
rect 5823 24157 5857 24191
rect 6929 24157 6963 24191
rect 7113 24157 7147 24191
rect 7849 24157 7883 24191
rect 8953 24157 8987 24191
rect 9227 24157 9261 24191
rect 10793 24157 10827 24191
rect 10977 24157 11011 24191
rect 1501 24089 1535 24123
rect 1685 24089 1719 24123
rect 13185 24089 13219 24123
rect 13553 24089 13587 24123
rect 6561 24021 6595 24055
rect 8769 24021 8803 24055
rect 8217 23817 8251 23851
rect 14473 23749 14507 23783
rect 4905 23681 4939 23715
rect 5179 23681 5213 23715
rect 6561 23681 6595 23715
rect 7297 23681 7331 23715
rect 7573 23681 7607 23715
rect 9379 23681 9413 23715
rect 12173 23681 12207 23715
rect 12633 23681 12667 23715
rect 13829 23681 13863 23715
rect 6377 23613 6411 23647
rect 7414 23613 7448 23647
rect 9137 23613 9171 23647
rect 12817 23613 12851 23647
rect 13553 23613 13587 23647
rect 13670 23613 13704 23647
rect 5917 23545 5951 23579
rect 7021 23545 7055 23579
rect 13277 23545 13311 23579
rect 10149 23477 10183 23511
rect 12449 23477 12483 23511
rect 11989 23273 12023 23307
rect 13369 23273 13403 23307
rect 10977 23137 11011 23171
rect 12357 23137 12391 23171
rect 1685 23069 1719 23103
rect 11251 23069 11285 23103
rect 12631 23069 12665 23103
rect 14197 23069 14231 23103
rect 1501 23001 1535 23035
rect 14381 22933 14415 22967
rect 1593 22729 1627 22763
rect 13369 22729 13403 22763
rect 14381 22729 14415 22763
rect 1501 22593 1535 22627
rect 8399 22593 8433 22627
rect 10057 22593 10091 22627
rect 10315 22623 10349 22657
rect 11713 22593 11747 22627
rect 12449 22593 12483 22627
rect 12587 22593 12621 22627
rect 12725 22593 12759 22627
rect 13553 22593 13587 22627
rect 14105 22593 14139 22627
rect 8125 22525 8159 22559
rect 11529 22525 11563 22559
rect 11069 22457 11103 22491
rect 12173 22457 12207 22491
rect 9137 22389 9171 22423
rect 13829 22389 13863 22423
rect 14289 22185 14323 22219
rect 7389 22049 7423 22083
rect 9781 22049 9815 22083
rect 10425 22049 10459 22083
rect 10701 22049 10735 22083
rect 10977 22049 11011 22083
rect 6009 21981 6043 22015
rect 6251 21981 6285 22015
rect 7663 21981 7697 22015
rect 9965 21981 9999 22015
rect 10839 21981 10873 22015
rect 12173 21981 12207 22015
rect 12431 21951 12465 21985
rect 14105 21981 14139 22015
rect 7021 21845 7055 21879
rect 8401 21845 8435 21879
rect 11621 21845 11655 21879
rect 13185 21845 13219 21879
rect 9873 21641 9907 21675
rect 11897 21641 11931 21675
rect 12541 21573 12575 21607
rect 1501 21505 1535 21539
rect 6635 21535 6669 21569
rect 8217 21505 8251 21539
rect 9229 21505 9263 21539
rect 11621 21505 11655 21539
rect 12173 21505 12207 21539
rect 13553 21505 13587 21539
rect 6377 21437 6411 21471
rect 8033 21437 8067 21471
rect 8677 21437 8711 21471
rect 8953 21437 8987 21471
rect 9091 21437 9125 21471
rect 12633 21437 12667 21471
rect 12817 21437 12851 21471
rect 13277 21437 13311 21471
rect 13670 21437 13704 21471
rect 13829 21437 13863 21471
rect 1685 21369 1719 21403
rect 7389 21301 7423 21335
rect 14473 21301 14507 21335
rect 3341 21097 3375 21131
rect 8217 21097 8251 21131
rect 11897 21097 11931 21131
rect 13645 21097 13679 21131
rect 1685 20961 1719 20995
rect 7021 20961 7055 20995
rect 7297 20961 7331 20995
rect 12633 20961 12667 20995
rect 1409 20893 1443 20927
rect 3157 20893 3191 20927
rect 6377 20893 6411 20927
rect 6561 20893 6595 20927
rect 7414 20893 7448 20927
rect 7573 20893 7607 20927
rect 9781 20893 9815 20927
rect 10023 20893 10057 20927
rect 11437 20893 11471 20927
rect 11621 20893 11655 20927
rect 12891 20893 12925 20927
rect 12173 20825 12207 20859
rect 12541 20825 12575 20859
rect 10793 20757 10827 20791
rect 11253 20757 11287 20791
rect 7021 20553 7055 20587
rect 11989 20553 12023 20587
rect 14013 20553 14047 20587
rect 13737 20485 13771 20519
rect 5069 20417 5103 20451
rect 6469 20417 6503 20451
rect 7205 20417 7239 20451
rect 7297 20417 7331 20451
rect 7481 20417 7515 20451
rect 8491 20417 8525 20451
rect 9839 20417 9873 20451
rect 11161 20417 11195 20451
rect 11345 20417 11379 20451
rect 11713 20417 11747 20451
rect 12447 20417 12481 20451
rect 4813 20349 4847 20383
rect 6653 20349 6687 20383
rect 8217 20349 8251 20383
rect 9597 20349 9631 20383
rect 12173 20349 12207 20383
rect 6193 20281 6227 20315
rect 7389 20213 7423 20247
rect 9229 20213 9263 20247
rect 10609 20213 10643 20247
rect 11253 20213 11287 20247
rect 13185 20213 13219 20247
rect 10793 20009 10827 20043
rect 11345 20009 11379 20043
rect 13921 20009 13955 20043
rect 1685 19941 1719 19975
rect 6837 19941 6871 19975
rect 8493 19941 8527 19975
rect 9597 19941 9631 19975
rect 12725 19941 12759 19975
rect 7481 19873 7515 19907
rect 8953 19873 8987 19907
rect 9873 19873 9907 19907
rect 10147 19873 10181 19907
rect 12081 19873 12115 19907
rect 13001 19873 13035 19907
rect 13139 19873 13173 19907
rect 5825 19805 5859 19839
rect 6099 19795 6133 19829
rect 7389 19805 7423 19839
rect 7723 19805 7757 19839
rect 9137 19805 9171 19839
rect 9990 19805 10024 19839
rect 11069 19805 11103 19839
rect 12265 19805 12299 19839
rect 13277 19805 13311 19839
rect 1501 19737 1535 19771
rect 11621 19737 11655 19771
rect 11989 19737 12023 19771
rect 7205 19669 7239 19703
rect 11069 19465 11103 19499
rect 13737 19465 13771 19499
rect 14381 19465 14415 19499
rect 7389 19397 7423 19431
rect 1501 19329 1535 19363
rect 6837 19329 6871 19363
rect 7021 19329 7055 19363
rect 7113 19329 7147 19363
rect 7481 19329 7515 19363
rect 8215 19329 8249 19363
rect 10793 19329 10827 19363
rect 11253 19329 11287 19363
rect 11529 19329 11563 19363
rect 12081 19329 12115 19363
rect 12725 19329 12759 19363
rect 12967 19329 13001 19363
rect 14197 19329 14231 19363
rect 6929 19261 6963 19295
rect 7392 19261 7426 19295
rect 7941 19261 7975 19295
rect 11805 19261 11839 19295
rect 1685 19193 1719 19227
rect 7205 19193 7239 19227
rect 7573 19193 7607 19227
rect 10885 19193 10919 19227
rect 11621 19193 11655 19227
rect 8953 19125 8987 19159
rect 11713 19125 11747 19159
rect 12357 19125 12391 19159
rect 5273 18921 5307 18955
rect 11897 18921 11931 18955
rect 12449 18921 12483 18955
rect 6469 18853 6503 18887
rect 7297 18853 7331 18887
rect 7113 18785 7147 18819
rect 12633 18785 12667 18819
rect 5457 18717 5491 18751
rect 5731 18717 5765 18751
rect 6837 18717 6871 18751
rect 6929 18717 6963 18751
rect 7481 18717 7515 18751
rect 7573 18717 7607 18751
rect 9873 18717 9907 18751
rect 10131 18687 10165 18721
rect 11437 18717 11471 18751
rect 12173 18717 12207 18751
rect 12875 18717 12909 18751
rect 14289 18717 14323 18751
rect 5181 18649 5215 18683
rect 7665 18649 7699 18683
rect 11621 18649 11655 18683
rect 7113 18581 7147 18615
rect 10885 18581 10919 18615
rect 11253 18581 11287 18615
rect 13645 18581 13679 18615
rect 14105 18581 14139 18615
rect 6837 18377 6871 18411
rect 11345 18377 11379 18411
rect 14473 18377 14507 18411
rect 1501 18241 1535 18275
rect 5069 18241 5103 18275
rect 7021 18241 7055 18275
rect 8827 18241 8861 18275
rect 11161 18241 11195 18275
rect 11529 18241 11563 18275
rect 11989 18241 12023 18275
rect 12173 18241 12207 18275
rect 12265 18241 12299 18275
rect 13829 18241 13863 18275
rect 4813 18173 4847 18207
rect 8585 18173 8619 18207
rect 11805 18173 11839 18207
rect 12081 18173 12115 18207
rect 12633 18173 12667 18207
rect 12817 18173 12851 18207
rect 13553 18173 13587 18207
rect 13670 18173 13704 18207
rect 1685 18105 1719 18139
rect 6193 18105 6227 18139
rect 11621 18105 11655 18139
rect 12357 18105 12391 18139
rect 13277 18105 13311 18139
rect 9597 18037 9631 18071
rect 11713 18037 11747 18071
rect 11621 17833 11655 17867
rect 11897 17833 11931 17867
rect 13277 17833 13311 17867
rect 13829 17833 13863 17867
rect 1685 17765 1719 17799
rect 11345 17765 11379 17799
rect 9413 17697 9447 17731
rect 6193 17629 6227 17663
rect 6451 17599 6485 17633
rect 9687 17629 9721 17663
rect 11161 17629 11195 17663
rect 11437 17629 11471 17663
rect 12265 17629 12299 17663
rect 12507 17629 12541 17663
rect 13645 17629 13679 17663
rect 1501 17561 1535 17595
rect 11805 17561 11839 17595
rect 7205 17493 7239 17527
rect 10425 17493 10459 17527
rect 1593 17289 1627 17323
rect 8953 17289 8987 17323
rect 11345 17289 11379 17323
rect 13277 17289 13311 17323
rect 13829 17289 13863 17323
rect 14381 17289 14415 17323
rect 14105 17221 14139 17255
rect 1501 17153 1535 17187
rect 7113 17153 7147 17187
rect 8171 17153 8205 17187
rect 9505 17153 9539 17187
rect 10425 17153 10459 17187
rect 10701 17153 10735 17187
rect 11863 17153 11897 17187
rect 13185 17153 13219 17187
rect 13553 17153 13587 17187
rect 7297 17085 7331 17119
rect 7757 17085 7791 17119
rect 8033 17085 8067 17119
rect 8309 17085 8343 17119
rect 9689 17085 9723 17119
rect 10563 17085 10597 17119
rect 11621 17085 11655 17119
rect 10149 17017 10183 17051
rect 12633 16949 12667 16983
rect 7757 16745 7791 16779
rect 11805 16745 11839 16779
rect 10609 16677 10643 16711
rect 13737 16677 13771 16711
rect 6745 16609 6779 16643
rect 9965 16609 9999 16643
rect 10885 16609 10919 16643
rect 11002 16609 11036 16643
rect 11897 16609 11931 16643
rect 12081 16609 12115 16643
rect 12541 16609 12575 16643
rect 1409 16541 1443 16575
rect 1683 16541 1717 16575
rect 7019 16541 7053 16575
rect 10149 16541 10183 16575
rect 11161 16541 11195 16575
rect 12817 16541 12851 16575
rect 12934 16541 12968 16575
rect 13093 16541 13127 16575
rect 14289 16541 14323 16575
rect 14473 16473 14507 16507
rect 2421 16405 2455 16439
rect 12541 16201 12575 16235
rect 14473 16201 14507 16235
rect 10425 16133 10459 16167
rect 1667 16095 1701 16129
rect 7447 16065 7481 16099
rect 8585 16065 8619 16099
rect 8769 16065 8803 16099
rect 11771 16065 11805 16099
rect 13151 16065 13185 16099
rect 14289 16065 14323 16099
rect 1409 15997 1443 16031
rect 7205 15997 7239 16031
rect 9505 15997 9539 16031
rect 9622 15997 9656 16031
rect 9781 15997 9815 16031
rect 11529 15997 11563 16031
rect 12909 15997 12943 16031
rect 8217 15929 8251 15963
rect 9229 15929 9263 15963
rect 2421 15861 2455 15895
rect 13921 15861 13955 15895
rect 1593 15657 1627 15691
rect 9965 15657 9999 15691
rect 14381 15657 14415 15691
rect 11989 15589 12023 15623
rect 12725 15589 12759 15623
rect 8953 15521 8987 15555
rect 12265 15521 12299 15555
rect 1501 15453 1535 15487
rect 1961 15453 1995 15487
rect 5457 15453 5491 15487
rect 5715 15443 5749 15477
rect 9227 15453 9261 15487
rect 10333 15453 10367 15487
rect 10591 15423 10625 15457
rect 11805 15453 11839 15487
rect 12081 15453 12115 15487
rect 13001 15453 13035 15487
rect 13118 15453 13152 15487
rect 13277 15453 13311 15487
rect 14289 15453 14323 15487
rect 13921 15385 13955 15419
rect 1777 15317 1811 15351
rect 6469 15317 6503 15351
rect 11345 15317 11379 15351
rect 6561 15113 6595 15147
rect 7665 15113 7699 15147
rect 7849 15113 7883 15147
rect 12817 15113 12851 15147
rect 14013 15113 14047 15147
rect 1501 15045 1535 15079
rect 6837 15045 6871 15079
rect 12725 15045 12759 15079
rect 2145 14977 2179 15011
rect 6929 14977 6963 15011
rect 7297 14977 7331 15011
rect 10023 14977 10057 15011
rect 11805 14977 11839 15011
rect 13243 14977 13277 15011
rect 9781 14909 9815 14943
rect 13001 14909 13035 14943
rect 11989 14841 12023 14875
rect 1593 14773 1627 14807
rect 1961 14773 1995 14807
rect 10793 14773 10827 14807
rect 6837 14569 6871 14603
rect 12265 14569 12299 14603
rect 14381 14569 14415 14603
rect 11069 14501 11103 14535
rect 5825 14433 5859 14467
rect 10425 14433 10459 14467
rect 10609 14433 10643 14467
rect 11462 14433 11496 14467
rect 11621 14433 11655 14467
rect 12633 14433 12667 14467
rect 1409 14365 1443 14399
rect 1683 14365 1717 14399
rect 6067 14365 6101 14399
rect 7205 14365 7239 14399
rect 7479 14365 7513 14399
rect 11345 14365 11379 14399
rect 12875 14365 12909 14399
rect 14289 14365 14323 14399
rect 2421 14229 2455 14263
rect 8217 14229 8251 14263
rect 13645 14229 13679 14263
rect 1593 14025 1627 14059
rect 8769 14025 8803 14059
rect 10333 14025 10367 14059
rect 14473 14025 14507 14059
rect 1501 13957 1535 13991
rect 9045 13957 9079 13991
rect 10149 13957 10183 13991
rect 2145 13889 2179 13923
rect 6929 13889 6963 13923
rect 8125 13889 8159 13923
rect 9321 13889 9355 13923
rect 9413 13889 9447 13923
rect 9781 13889 9815 13923
rect 11529 13889 11563 13923
rect 11803 13889 11837 13923
rect 13151 13889 13185 13923
rect 14289 13889 14323 13923
rect 7113 13821 7147 13855
rect 7849 13821 7883 13855
rect 7987 13821 8021 13855
rect 12909 13821 12943 13855
rect 7573 13753 7607 13787
rect 1961 13685 1995 13719
rect 12541 13685 12575 13719
rect 13921 13685 13955 13719
rect 7113 13481 7147 13515
rect 8493 13481 8527 13515
rect 9965 13481 9999 13515
rect 13369 13481 13403 13515
rect 13921 13481 13955 13515
rect 14381 13481 14415 13515
rect 12173 13413 12207 13447
rect 6101 13345 6135 13379
rect 7481 13345 7515 13379
rect 11713 13345 11747 13379
rect 12449 13345 12483 13379
rect 12587 13345 12621 13379
rect 1501 13277 1535 13311
rect 6359 13247 6393 13281
rect 7755 13277 7789 13311
rect 8953 13277 8987 13311
rect 9227 13277 9261 13311
rect 11529 13277 11563 13311
rect 12725 13277 12759 13311
rect 13461 13277 13495 13311
rect 13737 13277 13771 13311
rect 14289 13277 14323 13311
rect 1593 13141 1627 13175
rect 13645 13141 13679 13175
rect 11989 12937 12023 12971
rect 1683 12811 1717 12845
rect 11805 12801 11839 12835
rect 12081 12801 12115 12835
rect 12357 12801 12391 12835
rect 12817 12801 12851 12835
rect 13553 12801 13587 12835
rect 13829 12801 13863 12835
rect 1409 12733 1443 12767
rect 12633 12733 12667 12767
rect 13670 12733 13704 12767
rect 13277 12665 13311 12699
rect 14473 12665 14507 12699
rect 2421 12597 2455 12631
rect 12265 12597 12299 12631
rect 12541 12597 12575 12631
rect 1593 12393 1627 12427
rect 12449 12393 12483 12427
rect 13921 12393 13955 12427
rect 6561 12257 6595 12291
rect 11437 12257 11471 12291
rect 12817 12257 12851 12291
rect 2145 12189 2179 12223
rect 6803 12189 6837 12223
rect 11711 12189 11745 12223
rect 13093 12189 13127 12223
rect 13737 12189 13771 12223
rect 14289 12189 14323 12223
rect 1501 12121 1535 12155
rect 1961 12053 1995 12087
rect 7573 12053 7607 12087
rect 14473 12053 14507 12087
rect 10425 11849 10459 11883
rect 14473 11849 14507 11883
rect 9137 11781 9171 11815
rect 9505 11781 9539 11815
rect 10241 11781 10275 11815
rect 1501 11713 1535 11747
rect 5163 11743 5197 11777
rect 6929 11713 6963 11747
rect 7847 11713 7881 11747
rect 9413 11713 9447 11747
rect 9873 11713 9907 11747
rect 11989 11713 12023 11747
rect 13670 11713 13704 11747
rect 13829 11713 13863 11747
rect 4905 11645 4939 11679
rect 7573 11645 7607 11679
rect 11713 11645 11747 11679
rect 12633 11645 12667 11679
rect 12817 11645 12851 11679
rect 13553 11645 13587 11679
rect 8585 11577 8619 11611
rect 13277 11577 13311 11611
rect 1593 11509 1627 11543
rect 5917 11509 5951 11543
rect 7021 11509 7055 11543
rect 10057 11305 10091 11339
rect 13093 11305 13127 11339
rect 13921 11305 13955 11339
rect 14473 11305 14507 11339
rect 13645 11237 13679 11271
rect 5273 11169 5307 11203
rect 7573 11169 7607 11203
rect 7987 11169 8021 11203
rect 9045 11169 9079 11203
rect 11437 11169 11471 11203
rect 5547 11101 5581 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 7849 11101 7883 11135
rect 8125 11101 8159 11135
rect 9319 11101 9353 11135
rect 10885 11101 10919 11135
rect 11161 11101 11195 11135
rect 12081 11101 12115 11135
rect 12323 11101 12357 11135
rect 13461 11101 13495 11135
rect 13737 11101 13771 11135
rect 14289 11101 14323 11135
rect 1501 11033 1535 11067
rect 1593 10965 1627 10999
rect 6285 10965 6319 10999
rect 6653 10965 6687 10999
rect 8769 10965 8803 10999
rect 11069 10965 11103 10999
rect 1593 10761 1627 10795
rect 13829 10761 13863 10795
rect 14381 10761 14415 10795
rect 1777 10625 1811 10659
rect 5917 10625 5951 10659
rect 6561 10625 6595 10659
rect 7757 10625 7791 10659
rect 12449 10625 12483 10659
rect 13059 10625 13093 10659
rect 14197 10625 14231 10659
rect 6009 10557 6043 10591
rect 6193 10557 6227 10591
rect 6745 10557 6779 10591
rect 7481 10557 7515 10591
rect 7619 10557 7653 10591
rect 8677 10557 8711 10591
rect 11529 10557 11563 10591
rect 11805 10557 11839 10591
rect 12817 10557 12851 10591
rect 7205 10489 7239 10523
rect 6101 10421 6135 10455
rect 8401 10421 8435 10455
rect 12633 10421 12667 10455
rect 2421 10217 2455 10251
rect 6837 10217 6871 10251
rect 7849 10217 7883 10251
rect 11989 10217 12023 10251
rect 13921 10217 13955 10251
rect 2237 10149 2271 10183
rect 7573 10149 7607 10183
rect 14473 10149 14507 10183
rect 10057 10081 10091 10115
rect 10517 10081 10551 10115
rect 10910 10081 10944 10115
rect 11069 10081 11103 10115
rect 12081 10081 12115 10115
rect 12725 10081 12759 10115
rect 13001 10081 13035 10115
rect 13139 10081 13173 10115
rect 2053 10013 2087 10047
rect 2329 10013 2363 10047
rect 6745 10013 6779 10047
rect 6929 10013 6963 10047
rect 7757 10013 7791 10047
rect 8033 10013 8067 10047
rect 9873 10013 9907 10047
rect 10793 10013 10827 10047
rect 11805 10013 11839 10047
rect 12265 10013 12299 10047
rect 13277 10013 13311 10047
rect 1501 9945 1535 9979
rect 14289 9945 14323 9979
rect 1593 9877 1627 9911
rect 11713 9877 11747 9911
rect 2789 9673 2823 9707
rect 1683 9537 1717 9571
rect 2973 9537 3007 9571
rect 6469 9537 6503 9571
rect 6653 9537 6687 9571
rect 9505 9537 9539 9571
rect 9689 9537 9723 9571
rect 10425 9537 10459 9571
rect 10563 9537 10597 9571
rect 11713 9537 11747 9571
rect 12587 9537 12621 9571
rect 12725 9537 12759 9571
rect 13921 9537 13955 9571
rect 1409 9469 1443 9503
rect 8401 9469 8435 9503
rect 10701 9469 10735 9503
rect 11529 9469 11563 9503
rect 12449 9469 12483 9503
rect 13645 9469 13679 9503
rect 2421 9401 2455 9435
rect 10149 9401 10183 9435
rect 12173 9401 12207 9435
rect 6561 9333 6595 9367
rect 11345 9333 11379 9367
rect 13369 9333 13403 9367
rect 6745 9129 6779 9163
rect 14381 9129 14415 9163
rect 6193 9061 6227 9095
rect 11805 9061 11839 9095
rect 13921 9061 13955 9095
rect 5181 8993 5215 9027
rect 6837 8993 6871 9027
rect 6929 8993 6963 9027
rect 7573 8993 7607 9027
rect 7849 8993 7883 9027
rect 7987 8993 8021 9027
rect 8125 8993 8159 9027
rect 9873 8993 9907 9027
rect 10287 8993 10321 9027
rect 10425 8993 10459 9027
rect 12081 8993 12115 9027
rect 12219 8993 12253 9027
rect 1409 8925 1443 8959
rect 1667 8895 1701 8929
rect 5439 8895 5473 8929
rect 6561 8925 6595 8959
rect 6653 8925 6687 8959
rect 7113 8925 7147 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 9413 8925 9447 8959
rect 10167 8925 10201 8959
rect 11069 8925 11103 8959
rect 11161 8925 11195 8959
rect 11345 8925 11379 8959
rect 12357 8925 12391 8959
rect 13001 8925 13035 8959
rect 14289 8925 14323 8959
rect 13369 8857 13403 8891
rect 13737 8857 13771 8891
rect 2421 8789 2455 8823
rect 8769 8789 8803 8823
rect 13461 8789 13495 8823
rect 1961 8585 1995 8619
rect 6009 8585 6043 8619
rect 6561 8585 6595 8619
rect 6929 8585 6963 8619
rect 9229 8585 9263 8619
rect 12541 8585 12575 8619
rect 13921 8585 13955 8619
rect 1501 8517 1535 8551
rect 2145 8449 2179 8483
rect 6193 8449 6227 8483
rect 6469 8449 6503 8483
rect 7113 8449 7147 8483
rect 8309 8449 8343 8483
rect 9505 8449 9539 8483
rect 9689 8449 9723 8483
rect 10542 8449 10576 8483
rect 10701 8449 10735 8483
rect 11803 8449 11837 8483
rect 13167 8479 13201 8513
rect 7389 8381 7423 8415
rect 7573 8381 7607 8415
rect 8447 8381 8481 8415
rect 8595 8381 8629 8415
rect 10425 8381 10459 8415
rect 11529 8381 11563 8415
rect 12909 8381 12943 8415
rect 1685 8313 1719 8347
rect 8033 8313 8067 8347
rect 10149 8313 10183 8347
rect 11345 8313 11379 8347
rect 7849 8041 7883 8075
rect 12633 8041 12667 8075
rect 13829 8041 13863 8075
rect 14473 7973 14507 8007
rect 6837 7905 6871 7939
rect 10701 7905 10735 7939
rect 7095 7807 7129 7841
rect 10977 7837 11011 7871
rect 11621 7837 11655 7871
rect 11895 7837 11929 7871
rect 14289 7837 14323 7871
rect 1501 7769 1535 7803
rect 13737 7769 13771 7803
rect 1593 7701 1627 7735
rect 8769 7497 8803 7531
rect 11345 7497 11379 7531
rect 12541 7497 12575 7531
rect 14381 7497 14415 7531
rect 13093 7429 13127 7463
rect 13369 7429 13403 7463
rect 14197 7429 14231 7463
rect 1683 7361 1717 7395
rect 7999 7361 8033 7395
rect 9505 7361 9539 7395
rect 10701 7361 10735 7395
rect 11803 7361 11837 7395
rect 13461 7361 13495 7395
rect 13829 7361 13863 7395
rect 1409 7293 1443 7327
rect 7757 7293 7791 7327
rect 9689 7293 9723 7327
rect 10149 7293 10183 7327
rect 10425 7293 10459 7327
rect 10563 7293 10597 7327
rect 11529 7293 11563 7327
rect 2421 7157 2455 7191
rect 2421 6953 2455 6987
rect 13829 6885 13863 6919
rect 9413 6817 9447 6851
rect 9873 6817 9907 6851
rect 10149 6817 10183 6851
rect 10287 6817 10321 6851
rect 10425 6817 10459 6851
rect 11713 6817 11747 6851
rect 2329 6749 2363 6783
rect 2605 6749 2639 6783
rect 9229 6749 9263 6783
rect 11437 6749 11471 6783
rect 12817 6749 12851 6783
rect 12909 6749 12943 6783
rect 1501 6681 1535 6715
rect 13277 6681 13311 6715
rect 13645 6681 13679 6715
rect 14289 6681 14323 6715
rect 1593 6613 1627 6647
rect 2145 6613 2179 6647
rect 11069 6613 11103 6647
rect 12541 6613 12575 6647
rect 14381 6613 14415 6647
rect 2421 6409 2455 6443
rect 9137 6409 9171 6443
rect 1409 6273 1443 6307
rect 1683 6273 1717 6307
rect 8367 6273 8401 6307
rect 9505 6273 9539 6307
rect 10701 6273 10735 6307
rect 11529 6273 11563 6307
rect 12449 6273 12483 6307
rect 12566 6273 12600 6307
rect 12725 6273 12759 6307
rect 13645 6273 13679 6307
rect 8125 6205 8159 6239
rect 9689 6205 9723 6239
rect 10149 6205 10183 6239
rect 10425 6205 10459 6239
rect 10563 6205 10597 6239
rect 11345 6205 11379 6239
rect 11713 6205 11747 6239
rect 13921 6205 13955 6239
rect 12173 6137 12207 6171
rect 13369 6069 13403 6103
rect 1593 5865 1627 5899
rect 8493 5865 8527 5899
rect 11897 5865 11931 5899
rect 13277 5865 13311 5899
rect 13921 5797 13955 5831
rect 10885 5729 10919 5763
rect 12265 5729 12299 5763
rect 2053 5661 2087 5695
rect 2513 5661 2547 5695
rect 7481 5661 7515 5695
rect 7755 5661 7789 5695
rect 11127 5661 11161 5695
rect 12507 5661 12541 5695
rect 1501 5593 1535 5627
rect 13737 5593 13771 5627
rect 14289 5593 14323 5627
rect 2145 5525 2179 5559
rect 2329 5525 2363 5559
rect 14381 5525 14415 5559
rect 9137 5321 9171 5355
rect 10517 5321 10551 5355
rect 13369 5321 13403 5355
rect 1501 5253 1535 5287
rect 8125 5185 8159 5219
rect 8399 5185 8433 5219
rect 9779 5185 9813 5219
rect 12357 5185 12391 5219
rect 12631 5195 12665 5229
rect 9505 5117 9539 5151
rect 1593 4981 1627 5015
rect 1593 4777 1627 4811
rect 11621 4777 11655 4811
rect 13645 4777 13679 4811
rect 10609 4641 10643 4675
rect 1409 4573 1443 4607
rect 10851 4573 10885 4607
rect 12633 4573 12667 4607
rect 12875 4573 12909 4607
rect 13151 4097 13185 4131
rect 12909 4029 12943 4063
rect 13921 3893 13955 3927
rect 14289 3689 14323 3723
rect 13093 3553 13127 3587
rect 13369 3485 13403 3519
rect 14197 3485 14231 3519
rect 13645 3009 13679 3043
rect 13921 3009 13955 3043
rect 5825 2057 5859 2091
rect 6561 2057 6595 2091
rect 7297 2057 7331 2091
rect 8033 2057 8067 2091
rect 9413 2057 9447 2091
rect 10241 2057 10275 2091
rect 11713 2057 11747 2091
rect 12449 2057 12483 2091
rect 14197 2057 14231 2091
rect 8769 1989 8803 2023
rect 11069 1989 11103 2023
rect 14105 1989 14139 2023
rect 1409 1921 1443 1955
rect 3065 1921 3099 1955
rect 5733 1921 5767 1955
rect 6469 1921 6503 1955
rect 7205 1921 7239 1955
rect 7941 1921 7975 1955
rect 8585 1921 8619 1955
rect 9321 1921 9355 1955
rect 10149 1921 10183 1955
rect 10885 1921 10919 1955
rect 11621 1921 11655 1955
rect 12357 1921 12391 1955
rect 13001 1921 13035 1955
rect 13737 1921 13771 1955
rect 2237 1853 2271 1887
rect 3709 1853 3743 1887
rect 13921 1853 13955 1887
rect 13185 1785 13219 1819
rect 5825 1513 5859 1547
rect 6561 1513 6595 1547
rect 7297 1513 7331 1547
rect 8033 1513 8067 1547
rect 8953 1513 8987 1547
rect 9505 1513 9539 1547
rect 10241 1513 10275 1547
rect 10977 1513 11011 1547
rect 11713 1513 11747 1547
rect 12449 1513 12483 1547
rect 13185 1513 13219 1547
rect 13461 1513 13495 1547
rect 13737 1513 13771 1547
rect 12909 1445 12943 1479
rect 2973 1377 3007 1411
rect 2145 1309 2179 1343
rect 3801 1309 3835 1343
rect 4629 1309 4663 1343
rect 5365 1309 5399 1343
rect 6009 1309 6043 1343
rect 6745 1309 6779 1343
rect 7481 1309 7515 1343
rect 8217 1309 8251 1343
rect 9137 1309 9171 1343
rect 9689 1309 9723 1343
rect 10425 1309 10459 1343
rect 11161 1309 11195 1343
rect 11897 1309 11931 1343
rect 12633 1309 12667 1343
rect 13093 1309 13127 1343
rect 13369 1309 13403 1343
rect 13645 1309 13679 1343
rect 13921 1309 13955 1343
rect 4077 1241 4111 1275
rect 4445 1241 4479 1275
rect 5181 1241 5215 1275
rect 14197 1241 14231 1275
rect 14381 1241 14415 1275
<< metal1 >>
rect 1104 43546 14971 43568
rect 1104 43494 4376 43546
rect 4428 43494 4440 43546
rect 4492 43494 4504 43546
rect 4556 43494 4568 43546
rect 4620 43494 4632 43546
rect 4684 43494 7803 43546
rect 7855 43494 7867 43546
rect 7919 43494 7931 43546
rect 7983 43494 7995 43546
rect 8047 43494 8059 43546
rect 8111 43494 11230 43546
rect 11282 43494 11294 43546
rect 11346 43494 11358 43546
rect 11410 43494 11422 43546
rect 11474 43494 11486 43546
rect 11538 43494 14657 43546
rect 14709 43494 14721 43546
rect 14773 43494 14785 43546
rect 14837 43494 14849 43546
rect 14901 43494 14913 43546
rect 14965 43494 14971 43546
rect 1104 43472 14971 43494
rect 1578 43392 1584 43444
rect 1636 43392 1642 43444
rect 2314 43392 2320 43444
rect 2372 43392 2378 43444
rect 2866 43392 2872 43444
rect 2924 43392 2930 43444
rect 3421 43435 3479 43441
rect 3421 43401 3433 43435
rect 3467 43401 3479 43435
rect 3421 43395 3479 43401
rect 842 43324 848 43376
rect 900 43364 906 43376
rect 3436 43364 3464 43395
rect 3510 43392 3516 43444
rect 3568 43432 3574 43444
rect 3973 43435 4031 43441
rect 3973 43432 3985 43435
rect 3568 43404 3985 43432
rect 3568 43392 3574 43404
rect 3973 43401 3985 43404
rect 4019 43401 4031 43435
rect 3973 43395 4031 43401
rect 4246 43392 4252 43444
rect 4304 43432 4310 43444
rect 4525 43435 4583 43441
rect 4525 43432 4537 43435
rect 4304 43404 4537 43432
rect 4304 43392 4310 43404
rect 4525 43401 4537 43404
rect 4571 43401 4583 43435
rect 4525 43395 4583 43401
rect 5258 43392 5264 43444
rect 5316 43392 5322 43444
rect 5902 43392 5908 43444
rect 5960 43392 5966 43444
rect 6730 43392 6736 43444
rect 6788 43392 6794 43444
rect 7466 43392 7472 43444
rect 7524 43392 7530 43444
rect 8202 43392 8208 43444
rect 8260 43392 8266 43444
rect 8662 43392 8668 43444
rect 8720 43432 8726 43444
rect 9125 43435 9183 43441
rect 9125 43432 9137 43435
rect 8720 43404 9137 43432
rect 8720 43392 8726 43404
rect 9125 43401 9137 43404
rect 9171 43401 9183 43435
rect 9125 43395 9183 43401
rect 9398 43392 9404 43444
rect 9456 43432 9462 43444
rect 9677 43435 9735 43441
rect 9677 43432 9689 43435
rect 9456 43404 9689 43432
rect 9456 43392 9462 43404
rect 9677 43401 9689 43404
rect 9723 43401 9735 43435
rect 9677 43395 9735 43401
rect 10410 43392 10416 43444
rect 10468 43392 10474 43444
rect 10870 43392 10876 43444
rect 10928 43432 10934 43444
rect 11701 43435 11759 43441
rect 11701 43432 11713 43435
rect 10928 43404 11713 43432
rect 10928 43392 10934 43404
rect 11701 43401 11713 43404
rect 11747 43401 11759 43435
rect 11701 43395 11759 43401
rect 11882 43392 11888 43444
rect 11940 43432 11946 43444
rect 12253 43435 12311 43441
rect 12253 43432 12265 43435
rect 11940 43404 12265 43432
rect 11940 43392 11946 43404
rect 12253 43401 12265 43404
rect 12299 43401 12311 43435
rect 12253 43395 12311 43401
rect 12342 43392 12348 43444
rect 12400 43432 12406 43444
rect 12621 43435 12679 43441
rect 12621 43432 12633 43435
rect 12400 43404 12633 43432
rect 12400 43392 12406 43404
rect 12621 43401 12633 43404
rect 12667 43401 12679 43435
rect 12621 43395 12679 43401
rect 13078 43392 13084 43444
rect 13136 43432 13142 43444
rect 13265 43435 13323 43441
rect 13265 43432 13277 43435
rect 13136 43404 13277 43432
rect 13136 43392 13142 43404
rect 13265 43401 13277 43404
rect 13311 43401 13323 43435
rect 13265 43395 13323 43401
rect 13817 43435 13875 43441
rect 13817 43401 13829 43435
rect 13863 43432 13875 43435
rect 15286 43432 15292 43444
rect 13863 43404 15292 43432
rect 13863 43401 13875 43404
rect 13817 43395 13875 43401
rect 15286 43392 15292 43404
rect 15344 43392 15350 43444
rect 900 43336 3464 43364
rect 900 43324 906 43336
rect 1489 43299 1547 43305
rect 1489 43265 1501 43299
rect 1535 43296 1547 43299
rect 1762 43296 1768 43308
rect 1535 43268 1768 43296
rect 1535 43265 1547 43268
rect 1489 43259 1547 43265
rect 1762 43256 1768 43268
rect 1820 43256 1826 43308
rect 2130 43256 2136 43308
rect 2188 43256 2194 43308
rect 2777 43299 2835 43305
rect 2777 43265 2789 43299
rect 2823 43296 2835 43299
rect 3050 43296 3056 43308
rect 2823 43268 3056 43296
rect 2823 43265 2835 43268
rect 2777 43259 2835 43265
rect 3050 43256 3056 43268
rect 3108 43256 3114 43308
rect 3234 43256 3240 43308
rect 3292 43256 3298 43308
rect 3786 43256 3792 43308
rect 3844 43256 3850 43308
rect 4430 43256 4436 43308
rect 4488 43256 4494 43308
rect 5074 43256 5080 43308
rect 5132 43256 5138 43308
rect 5810 43256 5816 43308
rect 5868 43256 5874 43308
rect 6638 43256 6644 43308
rect 6696 43256 6702 43308
rect 7282 43256 7288 43308
rect 7340 43256 7346 43308
rect 8110 43256 8116 43308
rect 8168 43256 8174 43308
rect 8938 43256 8944 43308
rect 8996 43256 9002 43308
rect 9214 43256 9220 43308
rect 9272 43296 9278 43308
rect 9585 43299 9643 43305
rect 9585 43296 9597 43299
rect 9272 43268 9597 43296
rect 9272 43256 9278 43268
rect 9585 43265 9597 43268
rect 9631 43265 9643 43299
rect 9585 43259 9643 43265
rect 10226 43256 10232 43308
rect 10284 43256 10290 43308
rect 11606 43256 11612 43308
rect 11664 43256 11670 43308
rect 12066 43256 12072 43308
rect 12124 43256 12130 43308
rect 12526 43256 12532 43308
rect 12584 43256 12590 43308
rect 12802 43256 12808 43308
rect 12860 43296 12866 43308
rect 13081 43299 13139 43305
rect 13081 43296 13093 43299
rect 12860 43268 13093 43296
rect 12860 43256 12866 43268
rect 13081 43265 13093 43268
rect 13127 43265 13139 43299
rect 13081 43259 13139 43265
rect 13541 43299 13599 43305
rect 13541 43265 13553 43299
rect 13587 43296 13599 43299
rect 13722 43296 13728 43308
rect 13587 43268 13728 43296
rect 13587 43265 13599 43268
rect 13541 43259 13599 43265
rect 13722 43256 13728 43268
rect 13780 43256 13786 43308
rect 14277 43299 14335 43305
rect 14277 43265 14289 43299
rect 14323 43296 14335 43299
rect 15010 43296 15016 43308
rect 14323 43268 15016 43296
rect 14323 43265 14335 43268
rect 14277 43259 14335 43265
rect 15010 43256 15016 43268
rect 15068 43256 15074 43308
rect 14090 43052 14096 43104
rect 14148 43052 14154 43104
rect 1104 43002 14812 43024
rect 1104 42950 2663 43002
rect 2715 42950 2727 43002
rect 2779 42950 2791 43002
rect 2843 42950 2855 43002
rect 2907 42950 2919 43002
rect 2971 42950 6090 43002
rect 6142 42950 6154 43002
rect 6206 42950 6218 43002
rect 6270 42950 6282 43002
rect 6334 42950 6346 43002
rect 6398 42950 9517 43002
rect 9569 42950 9581 43002
rect 9633 42950 9645 43002
rect 9697 42950 9709 43002
rect 9761 42950 9773 43002
rect 9825 42950 12944 43002
rect 12996 42950 13008 43002
rect 13060 42950 13072 43002
rect 13124 42950 13136 43002
rect 13188 42950 13200 43002
rect 13252 42950 14812 43002
rect 1104 42928 14812 42950
rect 2869 42891 2927 42897
rect 2869 42857 2881 42891
rect 2915 42888 2927 42891
rect 3234 42888 3240 42900
rect 2915 42860 3240 42888
rect 2915 42857 2927 42860
rect 2869 42851 2927 42857
rect 3234 42848 3240 42860
rect 3292 42848 3298 42900
rect 3329 42891 3387 42897
rect 3329 42857 3341 42891
rect 3375 42888 3387 42891
rect 3786 42888 3792 42900
rect 3375 42860 3792 42888
rect 3375 42857 3387 42860
rect 3329 42851 3387 42857
rect 3786 42848 3792 42860
rect 3844 42848 3850 42900
rect 4157 42891 4215 42897
rect 4157 42857 4169 42891
rect 4203 42888 4215 42891
rect 4430 42888 4436 42900
rect 4203 42860 4436 42888
rect 4203 42857 4215 42860
rect 4157 42851 4215 42857
rect 4430 42848 4436 42860
rect 4488 42848 4494 42900
rect 4893 42891 4951 42897
rect 4893 42857 4905 42891
rect 4939 42888 4951 42891
rect 5074 42888 5080 42900
rect 4939 42860 5080 42888
rect 4939 42857 4951 42860
rect 4893 42851 4951 42857
rect 5074 42848 5080 42860
rect 5132 42848 5138 42900
rect 5629 42891 5687 42897
rect 5629 42857 5641 42891
rect 5675 42888 5687 42891
rect 5810 42888 5816 42900
rect 5675 42860 5816 42888
rect 5675 42857 5687 42860
rect 5629 42851 5687 42857
rect 5810 42848 5816 42860
rect 5868 42848 5874 42900
rect 6365 42891 6423 42897
rect 6365 42857 6377 42891
rect 6411 42888 6423 42891
rect 6638 42888 6644 42900
rect 6411 42860 6644 42888
rect 6411 42857 6423 42860
rect 6365 42851 6423 42857
rect 6638 42848 6644 42860
rect 6696 42848 6702 42900
rect 7101 42891 7159 42897
rect 7101 42857 7113 42891
rect 7147 42888 7159 42891
rect 7282 42888 7288 42900
rect 7147 42860 7288 42888
rect 7147 42857 7159 42860
rect 7101 42851 7159 42857
rect 7282 42848 7288 42860
rect 7340 42848 7346 42900
rect 7837 42891 7895 42897
rect 7837 42857 7849 42891
rect 7883 42888 7895 42891
rect 8110 42888 8116 42900
rect 7883 42860 8116 42888
rect 7883 42857 7895 42860
rect 7837 42851 7895 42857
rect 8110 42848 8116 42860
rect 8168 42848 8174 42900
rect 8573 42891 8631 42897
rect 8573 42857 8585 42891
rect 8619 42888 8631 42891
rect 8938 42888 8944 42900
rect 8619 42860 8944 42888
rect 8619 42857 8631 42860
rect 8573 42851 8631 42857
rect 8938 42848 8944 42860
rect 8996 42848 9002 42900
rect 9214 42848 9220 42900
rect 9272 42848 9278 42900
rect 10226 42848 10232 42900
rect 10284 42848 10290 42900
rect 10781 42891 10839 42897
rect 10781 42857 10793 42891
rect 10827 42888 10839 42891
rect 11606 42888 11612 42900
rect 10827 42860 11612 42888
rect 10827 42857 10839 42860
rect 10781 42851 10839 42857
rect 11606 42848 11612 42860
rect 11664 42848 11670 42900
rect 12066 42848 12072 42900
rect 12124 42848 12130 42900
rect 12253 42891 12311 42897
rect 12253 42857 12265 42891
rect 12299 42888 12311 42891
rect 12526 42888 12532 42900
rect 12299 42860 12532 42888
rect 12299 42857 12311 42860
rect 12253 42851 12311 42857
rect 12526 42848 12532 42860
rect 12584 42848 12590 42900
rect 12802 42848 12808 42900
rect 12860 42888 12866 42900
rect 12989 42891 13047 42897
rect 12989 42888 13001 42891
rect 12860 42860 13001 42888
rect 12860 42848 12866 42860
rect 12989 42857 13001 42860
rect 13035 42857 13047 42891
rect 12989 42851 13047 42857
rect 11517 42823 11575 42829
rect 11517 42789 11529 42823
rect 11563 42820 11575 42823
rect 12084 42820 12112 42848
rect 11563 42792 12112 42820
rect 11563 42789 11575 42792
rect 11517 42783 11575 42789
rect 3786 42712 3792 42764
rect 3844 42752 3850 42764
rect 13817 42755 13875 42761
rect 3844 42724 6592 42752
rect 3844 42712 3850 42724
rect 3510 42644 3516 42696
rect 3568 42644 3574 42696
rect 4062 42644 4068 42696
rect 4120 42684 4126 42696
rect 4341 42687 4399 42693
rect 4341 42684 4353 42687
rect 4120 42656 4353 42684
rect 4120 42644 4126 42656
rect 4341 42653 4353 42656
rect 4387 42653 4399 42687
rect 4341 42647 4399 42653
rect 5074 42644 5080 42696
rect 5132 42644 5138 42696
rect 6564 42693 6592 42724
rect 13817 42721 13829 42755
rect 13863 42752 13875 42755
rect 14550 42752 14556 42764
rect 13863 42724 14556 42752
rect 13863 42721 13875 42724
rect 13817 42715 13875 42721
rect 14550 42712 14556 42724
rect 14608 42712 14614 42764
rect 5813 42687 5871 42693
rect 5813 42653 5825 42687
rect 5859 42653 5871 42687
rect 5813 42647 5871 42653
rect 6549 42687 6607 42693
rect 6549 42653 6561 42687
rect 6595 42653 6607 42687
rect 6549 42647 6607 42653
rect 1397 42619 1455 42625
rect 1397 42585 1409 42619
rect 1443 42616 1455 42619
rect 4798 42616 4804 42628
rect 1443 42588 4804 42616
rect 1443 42585 1455 42588
rect 1397 42579 1455 42585
rect 4798 42576 4804 42588
rect 4856 42576 4862 42628
rect 3970 42508 3976 42560
rect 4028 42548 4034 42560
rect 5828 42548 5856 42647
rect 7282 42644 7288 42696
rect 7340 42644 7346 42696
rect 7466 42644 7472 42696
rect 7524 42684 7530 42696
rect 8021 42687 8079 42693
rect 8021 42684 8033 42687
rect 7524 42656 8033 42684
rect 7524 42644 7530 42656
rect 8021 42653 8033 42656
rect 8067 42653 8079 42687
rect 8021 42647 8079 42653
rect 8757 42687 8815 42693
rect 8757 42653 8769 42687
rect 8803 42653 8815 42687
rect 8757 42647 8815 42653
rect 7190 42576 7196 42628
rect 7248 42616 7254 42628
rect 8772 42616 8800 42647
rect 9398 42644 9404 42696
rect 9456 42644 9462 42696
rect 10045 42687 10103 42693
rect 10045 42684 10057 42687
rect 9692 42656 10057 42684
rect 7248 42588 8800 42616
rect 7248 42576 7254 42588
rect 4028 42520 5856 42548
rect 4028 42508 4034 42520
rect 8846 42508 8852 42560
rect 8904 42548 8910 42560
rect 9692 42557 9720 42656
rect 10045 42653 10057 42656
rect 10091 42653 10103 42687
rect 10045 42647 10103 42653
rect 10962 42644 10968 42696
rect 11020 42644 11026 42696
rect 11698 42644 11704 42696
rect 11756 42644 11762 42696
rect 12434 42644 12440 42696
rect 12492 42644 12498 42696
rect 13173 42687 13231 42693
rect 13173 42653 13185 42687
rect 13219 42684 13231 42687
rect 14277 42687 14335 42693
rect 13219 42656 13676 42684
rect 13219 42653 13231 42656
rect 13173 42647 13231 42653
rect 13538 42576 13544 42628
rect 13596 42576 13602 42628
rect 13648 42616 13676 42656
rect 14277 42653 14289 42687
rect 14323 42684 14335 42687
rect 15286 42684 15292 42696
rect 14323 42656 15292 42684
rect 14323 42653 14335 42656
rect 14277 42647 14335 42653
rect 15286 42644 15292 42656
rect 15344 42644 15350 42696
rect 15194 42616 15200 42628
rect 13648 42588 15200 42616
rect 15194 42576 15200 42588
rect 15252 42576 15258 42628
rect 9677 42551 9735 42557
rect 9677 42548 9689 42551
rect 8904 42520 9689 42548
rect 8904 42508 8910 42520
rect 9677 42517 9689 42520
rect 9723 42517 9735 42551
rect 9677 42511 9735 42517
rect 13722 42508 13728 42560
rect 13780 42548 13786 42560
rect 14093 42551 14151 42557
rect 14093 42548 14105 42551
rect 13780 42520 14105 42548
rect 13780 42508 13786 42520
rect 14093 42517 14105 42520
rect 14139 42517 14151 42551
rect 14093 42511 14151 42517
rect 1104 42458 14971 42480
rect 1104 42406 4376 42458
rect 4428 42406 4440 42458
rect 4492 42406 4504 42458
rect 4556 42406 4568 42458
rect 4620 42406 4632 42458
rect 4684 42406 7803 42458
rect 7855 42406 7867 42458
rect 7919 42406 7931 42458
rect 7983 42406 7995 42458
rect 8047 42406 8059 42458
rect 8111 42406 11230 42458
rect 11282 42406 11294 42458
rect 11346 42406 11358 42458
rect 11410 42406 11422 42458
rect 11474 42406 11486 42458
rect 11538 42406 14657 42458
rect 14709 42406 14721 42458
rect 14773 42406 14785 42458
rect 14837 42406 14849 42458
rect 14901 42406 14913 42458
rect 14965 42406 14971 42458
rect 1104 42384 14971 42406
rect 2041 42347 2099 42353
rect 2041 42313 2053 42347
rect 2087 42344 2099 42347
rect 2130 42344 2136 42356
rect 2087 42316 2136 42344
rect 2087 42313 2099 42316
rect 2041 42307 2099 42313
rect 2130 42304 2136 42316
rect 2188 42304 2194 42356
rect 4062 42304 4068 42356
rect 4120 42304 4126 42356
rect 4893 42347 4951 42353
rect 4893 42313 4905 42347
rect 4939 42344 4951 42347
rect 5074 42344 5080 42356
rect 4939 42316 5080 42344
rect 4939 42313 4951 42316
rect 4893 42307 4951 42313
rect 5074 42304 5080 42316
rect 5132 42304 5138 42356
rect 7190 42344 7196 42356
rect 6886 42316 7196 42344
rect 3878 42236 3884 42288
rect 3936 42276 3942 42288
rect 6886 42276 6914 42316
rect 7190 42304 7196 42316
rect 7248 42304 7254 42356
rect 7282 42304 7288 42356
rect 7340 42304 7346 42356
rect 7466 42304 7472 42356
rect 7524 42304 7530 42356
rect 13538 42304 13544 42356
rect 13596 42344 13602 42356
rect 13725 42347 13783 42353
rect 13725 42344 13737 42347
rect 13596 42316 13737 42344
rect 13596 42304 13602 42316
rect 13725 42313 13737 42316
rect 13771 42313 13783 42347
rect 13725 42307 13783 42313
rect 13814 42304 13820 42356
rect 13872 42344 13878 42356
rect 14185 42347 14243 42353
rect 14185 42344 14197 42347
rect 13872 42316 14197 42344
rect 13872 42304 13878 42316
rect 14185 42313 14197 42316
rect 14231 42313 14243 42347
rect 14185 42307 14243 42313
rect 3936 42248 6914 42276
rect 3936 42236 3942 42248
rect 2222 42168 2228 42220
rect 2280 42168 2286 42220
rect 4246 42168 4252 42220
rect 4304 42168 4310 42220
rect 5074 42168 5080 42220
rect 5132 42168 5138 42220
rect 4062 42100 4068 42152
rect 4120 42140 4126 42152
rect 7300 42140 7328 42304
rect 4120 42112 7328 42140
rect 4120 42100 4126 42112
rect 1026 42032 1032 42084
rect 1084 42072 1090 42084
rect 7484 42072 7512 42304
rect 14090 42236 14096 42288
rect 14148 42236 14154 42288
rect 13906 42168 13912 42220
rect 13964 42168 13970 42220
rect 1084 42044 7512 42072
rect 1084 42032 1090 42044
rect 1104 41914 14812 41936
rect 1104 41862 2663 41914
rect 2715 41862 2727 41914
rect 2779 41862 2791 41914
rect 2843 41862 2855 41914
rect 2907 41862 2919 41914
rect 2971 41862 6090 41914
rect 6142 41862 6154 41914
rect 6206 41862 6218 41914
rect 6270 41862 6282 41914
rect 6334 41862 6346 41914
rect 6398 41862 9517 41914
rect 9569 41862 9581 41914
rect 9633 41862 9645 41914
rect 9697 41862 9709 41914
rect 9761 41862 9773 41914
rect 9825 41862 12944 41914
rect 12996 41862 13008 41914
rect 13060 41862 13072 41914
rect 13124 41862 13136 41914
rect 13188 41862 13200 41914
rect 13252 41862 14812 41914
rect 1104 41840 14812 41862
rect 4154 41760 4160 41812
rect 4212 41800 4218 41812
rect 8846 41800 8852 41812
rect 4212 41772 8852 41800
rect 4212 41760 4218 41772
rect 8846 41760 8852 41772
rect 8904 41760 8910 41812
rect 1104 41370 14971 41392
rect 1104 41318 4376 41370
rect 4428 41318 4440 41370
rect 4492 41318 4504 41370
rect 4556 41318 4568 41370
rect 4620 41318 4632 41370
rect 4684 41318 7803 41370
rect 7855 41318 7867 41370
rect 7919 41318 7931 41370
rect 7983 41318 7995 41370
rect 8047 41318 8059 41370
rect 8111 41318 11230 41370
rect 11282 41318 11294 41370
rect 11346 41318 11358 41370
rect 11410 41318 11422 41370
rect 11474 41318 11486 41370
rect 11538 41318 14657 41370
rect 14709 41318 14721 41370
rect 14773 41318 14785 41370
rect 14837 41318 14849 41370
rect 14901 41318 14913 41370
rect 14965 41318 14971 41370
rect 1104 41296 14971 41318
rect 750 41080 756 41132
rect 808 41120 814 41132
rect 1397 41123 1455 41129
rect 1397 41120 1409 41123
rect 808 41092 1409 41120
rect 808 41080 814 41092
rect 1397 41089 1409 41092
rect 1443 41089 1455 41123
rect 1397 41083 1455 41089
rect 1581 40919 1639 40925
rect 1581 40885 1593 40919
rect 1627 40916 1639 40919
rect 9306 40916 9312 40928
rect 1627 40888 9312 40916
rect 1627 40885 1639 40888
rect 1581 40879 1639 40885
rect 9306 40876 9312 40888
rect 9364 40876 9370 40928
rect 1104 40826 14812 40848
rect 1104 40774 2663 40826
rect 2715 40774 2727 40826
rect 2779 40774 2791 40826
rect 2843 40774 2855 40826
rect 2907 40774 2919 40826
rect 2971 40774 6090 40826
rect 6142 40774 6154 40826
rect 6206 40774 6218 40826
rect 6270 40774 6282 40826
rect 6334 40774 6346 40826
rect 6398 40774 9517 40826
rect 9569 40774 9581 40826
rect 9633 40774 9645 40826
rect 9697 40774 9709 40826
rect 9761 40774 9773 40826
rect 9825 40774 12944 40826
rect 12996 40774 13008 40826
rect 13060 40774 13072 40826
rect 13124 40774 13136 40826
rect 13188 40774 13200 40826
rect 13252 40774 14812 40826
rect 1104 40752 14812 40774
rect 750 40468 756 40520
rect 808 40508 814 40520
rect 1397 40511 1455 40517
rect 1397 40508 1409 40511
rect 808 40480 1409 40508
rect 808 40468 814 40480
rect 1397 40477 1409 40480
rect 1443 40477 1455 40511
rect 1397 40471 1455 40477
rect 13538 40400 13544 40452
rect 13596 40400 13602 40452
rect 1581 40375 1639 40381
rect 1581 40341 1593 40375
rect 1627 40372 1639 40375
rect 5166 40372 5172 40384
rect 1627 40344 5172 40372
rect 1627 40341 1639 40344
rect 1581 40335 1639 40341
rect 5166 40332 5172 40344
rect 5224 40332 5230 40384
rect 13722 40332 13728 40384
rect 13780 40372 13786 40384
rect 13817 40375 13875 40381
rect 13817 40372 13829 40375
rect 13780 40344 13829 40372
rect 13780 40332 13786 40344
rect 13817 40341 13829 40344
rect 13863 40341 13875 40375
rect 13817 40335 13875 40341
rect 1104 40282 14971 40304
rect 1104 40230 4376 40282
rect 4428 40230 4440 40282
rect 4492 40230 4504 40282
rect 4556 40230 4568 40282
rect 4620 40230 4632 40282
rect 4684 40230 7803 40282
rect 7855 40230 7867 40282
rect 7919 40230 7931 40282
rect 7983 40230 7995 40282
rect 8047 40230 8059 40282
rect 8111 40230 11230 40282
rect 11282 40230 11294 40282
rect 11346 40230 11358 40282
rect 11410 40230 11422 40282
rect 11474 40230 11486 40282
rect 11538 40230 14657 40282
rect 14709 40230 14721 40282
rect 14773 40230 14785 40282
rect 14837 40230 14849 40282
rect 14901 40230 14913 40282
rect 14965 40230 14971 40282
rect 1104 40208 14971 40230
rect 9217 40171 9275 40177
rect 9217 40137 9229 40171
rect 9263 40137 9275 40171
rect 9217 40131 9275 40137
rect 10045 40171 10103 40177
rect 10045 40137 10057 40171
rect 10091 40168 10103 40171
rect 13538 40168 13544 40180
rect 10091 40140 13544 40168
rect 10091 40137 10103 40140
rect 10045 40131 10103 40137
rect 9232 40100 9260 40131
rect 13538 40128 13544 40140
rect 13596 40128 13602 40180
rect 9232 40072 10272 40100
rect 9306 39992 9312 40044
rect 9364 40032 9370 40044
rect 10244 40041 10272 40072
rect 9401 40035 9459 40041
rect 9401 40032 9413 40035
rect 9364 40004 9413 40032
rect 9364 39992 9370 40004
rect 9401 40001 9413 40004
rect 9447 40001 9459 40035
rect 9401 39995 9459 40001
rect 10229 40035 10287 40041
rect 10229 40001 10241 40035
rect 10275 40001 10287 40035
rect 10229 39995 10287 40001
rect 13354 39992 13360 40044
rect 13412 39992 13418 40044
rect 13906 39992 13912 40044
rect 13964 39992 13970 40044
rect 13633 39831 13691 39837
rect 13633 39797 13645 39831
rect 13679 39828 13691 39831
rect 13998 39828 14004 39840
rect 13679 39800 14004 39828
rect 13679 39797 13691 39800
rect 13633 39791 13691 39797
rect 13998 39788 14004 39800
rect 14056 39788 14062 39840
rect 14182 39788 14188 39840
rect 14240 39788 14246 39840
rect 1104 39738 14812 39760
rect 1104 39686 2663 39738
rect 2715 39686 2727 39738
rect 2779 39686 2791 39738
rect 2843 39686 2855 39738
rect 2907 39686 2919 39738
rect 2971 39686 6090 39738
rect 6142 39686 6154 39738
rect 6206 39686 6218 39738
rect 6270 39686 6282 39738
rect 6334 39686 6346 39738
rect 6398 39686 9517 39738
rect 9569 39686 9581 39738
rect 9633 39686 9645 39738
rect 9697 39686 9709 39738
rect 9761 39686 9773 39738
rect 9825 39686 12944 39738
rect 12996 39686 13008 39738
rect 13060 39686 13072 39738
rect 13124 39686 13136 39738
rect 13188 39686 13200 39738
rect 13252 39686 14812 39738
rect 1104 39664 14812 39686
rect 12989 39627 13047 39633
rect 12989 39593 13001 39627
rect 13035 39624 13047 39627
rect 13354 39624 13360 39636
rect 13035 39596 13360 39624
rect 13035 39593 13047 39596
rect 12989 39587 13047 39593
rect 13354 39584 13360 39596
rect 13412 39584 13418 39636
rect 8941 39559 8999 39565
rect 8941 39525 8953 39559
rect 8987 39525 8999 39559
rect 8941 39519 8999 39525
rect 9493 39559 9551 39565
rect 9493 39525 9505 39559
rect 9539 39556 9551 39559
rect 13906 39556 13912 39568
rect 9539 39528 13912 39556
rect 9539 39525 9551 39528
rect 9493 39519 9551 39525
rect 8956 39488 8984 39519
rect 13906 39516 13912 39528
rect 13964 39516 13970 39568
rect 8956 39460 9720 39488
rect 750 39380 756 39432
rect 808 39420 814 39432
rect 1397 39423 1455 39429
rect 1397 39420 1409 39423
rect 808 39392 1409 39420
rect 808 39380 814 39392
rect 1397 39389 1409 39392
rect 1443 39389 1455 39423
rect 1397 39383 1455 39389
rect 5166 39380 5172 39432
rect 5224 39420 5230 39432
rect 9692 39429 9720 39460
rect 9125 39423 9183 39429
rect 9125 39420 9137 39423
rect 5224 39392 9137 39420
rect 5224 39380 5230 39392
rect 9125 39389 9137 39392
rect 9171 39389 9183 39423
rect 9125 39383 9183 39389
rect 9677 39423 9735 39429
rect 9677 39389 9689 39423
rect 9723 39389 9735 39423
rect 9677 39383 9735 39389
rect 12802 39380 12808 39432
rect 12860 39420 12866 39432
rect 12897 39423 12955 39429
rect 12897 39420 12909 39423
rect 12860 39392 12909 39420
rect 12860 39380 12866 39392
rect 12897 39389 12909 39392
rect 12943 39389 12955 39423
rect 12897 39383 12955 39389
rect 13173 39423 13231 39429
rect 13173 39389 13185 39423
rect 13219 39389 13231 39423
rect 13173 39383 13231 39389
rect 13188 39352 13216 39383
rect 13262 39380 13268 39432
rect 13320 39420 13326 39432
rect 14185 39423 14243 39429
rect 14185 39420 14197 39423
rect 13320 39392 14197 39420
rect 13320 39380 13326 39392
rect 14185 39389 14197 39392
rect 14231 39389 14243 39423
rect 14185 39383 14243 39389
rect 12728 39324 13216 39352
rect 1578 39244 1584 39296
rect 1636 39244 1642 39296
rect 12728 39293 12756 39324
rect 13538 39312 13544 39364
rect 13596 39312 13602 39364
rect 13906 39312 13912 39364
rect 13964 39312 13970 39364
rect 12713 39287 12771 39293
rect 12713 39253 12725 39287
rect 12759 39253 12771 39287
rect 12713 39247 12771 39253
rect 14366 39244 14372 39296
rect 14424 39244 14430 39296
rect 1104 39194 14971 39216
rect 1104 39142 4376 39194
rect 4428 39142 4440 39194
rect 4492 39142 4504 39194
rect 4556 39142 4568 39194
rect 4620 39142 4632 39194
rect 4684 39142 7803 39194
rect 7855 39142 7867 39194
rect 7919 39142 7931 39194
rect 7983 39142 7995 39194
rect 8047 39142 8059 39194
rect 8111 39142 11230 39194
rect 11282 39142 11294 39194
rect 11346 39142 11358 39194
rect 11410 39142 11422 39194
rect 11474 39142 11486 39194
rect 11538 39142 14657 39194
rect 14709 39142 14721 39194
rect 14773 39142 14785 39194
rect 14837 39142 14849 39194
rect 14901 39142 14913 39194
rect 14965 39142 14971 39194
rect 1104 39120 14971 39142
rect 1578 39040 1584 39092
rect 1636 39080 1642 39092
rect 12713 39083 12771 39089
rect 1636 39052 2774 39080
rect 1636 39040 1642 39052
rect 2746 39012 2774 39052
rect 12713 39049 12725 39083
rect 12759 39080 12771 39083
rect 13538 39080 13544 39092
rect 12759 39052 13544 39080
rect 12759 39049 12771 39052
rect 12713 39043 12771 39049
rect 13538 39040 13544 39052
rect 13596 39040 13602 39092
rect 12802 39012 12808 39024
rect 2746 38984 12808 39012
rect 12802 38972 12808 38984
rect 12860 39012 12866 39024
rect 12860 38984 13584 39012
rect 12860 38972 12866 38984
rect 1394 38904 1400 38956
rect 1452 38904 1458 38956
rect 12710 38904 12716 38956
rect 12768 38944 12774 38956
rect 12897 38947 12955 38953
rect 12897 38944 12909 38947
rect 12768 38916 12909 38944
rect 12768 38904 12774 38916
rect 12897 38913 12909 38916
rect 12943 38913 12955 38947
rect 12897 38907 12955 38913
rect 13173 38947 13231 38953
rect 13173 38913 13185 38947
rect 13219 38913 13231 38947
rect 13173 38907 13231 38913
rect 12342 38836 12348 38888
rect 12400 38876 12406 38888
rect 13188 38876 13216 38907
rect 13354 38904 13360 38956
rect 13412 38904 13418 38956
rect 13556 38888 13584 38984
rect 13909 38947 13967 38953
rect 13909 38913 13921 38947
rect 13955 38944 13967 38947
rect 13998 38944 14004 38956
rect 13955 38916 14004 38944
rect 13955 38913 13967 38916
rect 13909 38907 13967 38913
rect 13998 38904 14004 38916
rect 14056 38904 14062 38956
rect 12400 38848 13216 38876
rect 12400 38836 12406 38848
rect 13538 38836 13544 38888
rect 13596 38836 13602 38888
rect 12989 38811 13047 38817
rect 12989 38777 13001 38811
rect 13035 38808 13047 38811
rect 13814 38808 13820 38820
rect 13035 38780 13820 38808
rect 13035 38777 13047 38780
rect 12989 38771 13047 38777
rect 13814 38768 13820 38780
rect 13872 38768 13878 38820
rect 1581 38743 1639 38749
rect 1581 38709 1593 38743
rect 1627 38740 1639 38743
rect 12802 38740 12808 38752
rect 1627 38712 12808 38740
rect 1627 38709 1639 38712
rect 1581 38703 1639 38709
rect 12802 38700 12808 38712
rect 12860 38700 12866 38752
rect 13630 38700 13636 38752
rect 13688 38700 13694 38752
rect 14182 38700 14188 38752
rect 14240 38700 14246 38752
rect 1104 38650 14812 38672
rect 1104 38598 2663 38650
rect 2715 38598 2727 38650
rect 2779 38598 2791 38650
rect 2843 38598 2855 38650
rect 2907 38598 2919 38650
rect 2971 38598 6090 38650
rect 6142 38598 6154 38650
rect 6206 38598 6218 38650
rect 6270 38598 6282 38650
rect 6334 38598 6346 38650
rect 6398 38598 9517 38650
rect 9569 38598 9581 38650
rect 9633 38598 9645 38650
rect 9697 38598 9709 38650
rect 9761 38598 9773 38650
rect 9825 38598 12944 38650
rect 12996 38598 13008 38650
rect 13060 38598 13072 38650
rect 13124 38598 13136 38650
rect 13188 38598 13200 38650
rect 13252 38598 14812 38650
rect 1104 38576 14812 38598
rect 12710 38496 12716 38548
rect 12768 38496 12774 38548
rect 13262 38496 13268 38548
rect 13320 38496 13326 38548
rect 12437 38471 12495 38477
rect 12437 38437 12449 38471
rect 12483 38468 12495 38471
rect 13280 38468 13308 38496
rect 12483 38440 13308 38468
rect 12483 38437 12495 38440
rect 12437 38431 12495 38437
rect 12710 38360 12716 38412
rect 12768 38400 12774 38412
rect 12768 38372 13216 38400
rect 12768 38360 12774 38372
rect 12618 38292 12624 38344
rect 12676 38292 12682 38344
rect 13188 38341 13216 38372
rect 12897 38335 12955 38341
rect 12897 38332 12909 38335
rect 12820 38304 12909 38332
rect 12820 38208 12848 38304
rect 12897 38301 12909 38304
rect 12943 38301 12955 38335
rect 12897 38295 12955 38301
rect 13173 38335 13231 38341
rect 13173 38301 13185 38335
rect 13219 38301 13231 38335
rect 13173 38295 13231 38301
rect 13446 38292 13452 38344
rect 13504 38292 13510 38344
rect 13633 38335 13691 38341
rect 13633 38301 13645 38335
rect 13679 38332 13691 38335
rect 13814 38332 13820 38344
rect 13679 38304 13820 38332
rect 13679 38301 13691 38304
rect 13633 38295 13691 38301
rect 13814 38292 13820 38304
rect 13872 38292 13878 38344
rect 14185 38335 14243 38341
rect 14185 38301 14197 38335
rect 14231 38301 14243 38335
rect 14185 38295 14243 38301
rect 14200 38264 14228 38295
rect 13004 38236 14228 38264
rect 12802 38156 12808 38208
rect 12860 38156 12866 38208
rect 13004 38205 13032 38236
rect 12989 38199 13047 38205
rect 12989 38165 13001 38199
rect 13035 38165 13047 38199
rect 12989 38159 13047 38165
rect 13262 38156 13268 38208
rect 13320 38156 13326 38208
rect 13814 38156 13820 38208
rect 13872 38156 13878 38208
rect 14366 38156 14372 38208
rect 14424 38156 14430 38208
rect 1104 38106 14971 38128
rect 1104 38054 4376 38106
rect 4428 38054 4440 38106
rect 4492 38054 4504 38106
rect 4556 38054 4568 38106
rect 4620 38054 4632 38106
rect 4684 38054 7803 38106
rect 7855 38054 7867 38106
rect 7919 38054 7931 38106
rect 7983 38054 7995 38106
rect 8047 38054 8059 38106
rect 8111 38054 11230 38106
rect 11282 38054 11294 38106
rect 11346 38054 11358 38106
rect 11410 38054 11422 38106
rect 11474 38054 11486 38106
rect 11538 38054 14657 38106
rect 14709 38054 14721 38106
rect 14773 38054 14785 38106
rect 14837 38054 14849 38106
rect 14901 38054 14913 38106
rect 14965 38054 14971 38106
rect 1104 38032 14971 38054
rect 11517 37995 11575 38001
rect 11517 37961 11529 37995
rect 11563 37961 11575 37995
rect 11517 37955 11575 37961
rect 11793 37995 11851 38001
rect 11793 37961 11805 37995
rect 11839 37992 11851 37995
rect 12618 37992 12624 38004
rect 11839 37964 12624 37992
rect 11839 37961 11851 37964
rect 11793 37955 11851 37961
rect 11532 37924 11560 37955
rect 12618 37952 12624 37964
rect 12676 37952 12682 38004
rect 12728 37964 14044 37992
rect 12728 37924 12756 37964
rect 14016 37936 14044 37964
rect 13262 37924 13268 37936
rect 11532 37896 12756 37924
rect 12820 37896 13268 37924
rect 750 37816 756 37868
rect 808 37856 814 37868
rect 1397 37859 1455 37865
rect 1397 37856 1409 37859
rect 808 37828 1409 37856
rect 808 37816 814 37828
rect 1397 37825 1409 37828
rect 1443 37825 1455 37859
rect 1397 37819 1455 37825
rect 10778 37816 10784 37868
rect 10836 37856 10842 37868
rect 12820 37865 12848 37896
rect 13262 37884 13268 37896
rect 13320 37884 13326 37936
rect 13998 37884 14004 37936
rect 14056 37884 14062 37936
rect 11701 37859 11759 37865
rect 11701 37856 11713 37859
rect 10836 37828 11713 37856
rect 10836 37816 10842 37828
rect 11701 37825 11713 37828
rect 11747 37825 11759 37859
rect 11701 37819 11759 37825
rect 11977 37859 12035 37865
rect 11977 37825 11989 37859
rect 12023 37825 12035 37859
rect 11977 37819 12035 37825
rect 12805 37859 12863 37865
rect 12805 37825 12817 37859
rect 12851 37825 12863 37859
rect 12805 37819 12863 37825
rect 12989 37859 13047 37865
rect 12989 37825 13001 37859
rect 13035 37825 13047 37859
rect 12989 37819 13047 37825
rect 13357 37859 13415 37865
rect 13357 37825 13369 37859
rect 13403 37825 13415 37859
rect 13357 37819 13415 37825
rect 1581 37723 1639 37729
rect 1581 37689 1593 37723
rect 1627 37720 1639 37723
rect 7650 37720 7656 37732
rect 1627 37692 7656 37720
rect 1627 37689 1639 37692
rect 1581 37683 1639 37689
rect 7650 37680 7656 37692
rect 7708 37720 7714 37732
rect 11992 37720 12020 37819
rect 12618 37748 12624 37800
rect 12676 37788 12682 37800
rect 13004 37788 13032 37819
rect 12676 37760 13032 37788
rect 13372 37788 13400 37819
rect 13538 37816 13544 37868
rect 13596 37816 13602 37868
rect 14093 37859 14151 37865
rect 14093 37825 14105 37859
rect 14139 37825 14151 37859
rect 14093 37819 14151 37825
rect 13998 37788 14004 37800
rect 13372 37760 14004 37788
rect 12676 37748 12682 37760
rect 13998 37748 14004 37760
rect 14056 37748 14062 37800
rect 7708 37692 12020 37720
rect 7708 37680 7714 37692
rect 12250 37680 12256 37732
rect 12308 37720 12314 37732
rect 14108 37720 14136 37819
rect 12308 37692 14136 37720
rect 12308 37680 12314 37692
rect 12621 37655 12679 37661
rect 12621 37621 12633 37655
rect 12667 37652 12679 37655
rect 13354 37652 13360 37664
rect 12667 37624 13360 37652
rect 12667 37621 12679 37624
rect 12621 37615 12679 37621
rect 13354 37612 13360 37624
rect 13412 37612 13418 37664
rect 13722 37612 13728 37664
rect 13780 37652 13786 37664
rect 13817 37655 13875 37661
rect 13817 37652 13829 37655
rect 13780 37624 13829 37652
rect 13780 37612 13786 37624
rect 13817 37621 13829 37624
rect 13863 37621 13875 37655
rect 13817 37615 13875 37621
rect 14369 37655 14427 37661
rect 14369 37621 14381 37655
rect 14415 37652 14427 37655
rect 15102 37652 15108 37664
rect 14415 37624 15108 37652
rect 14415 37621 14427 37624
rect 14369 37615 14427 37621
rect 15102 37612 15108 37624
rect 15160 37612 15166 37664
rect 1104 37562 14812 37584
rect 1104 37510 2663 37562
rect 2715 37510 2727 37562
rect 2779 37510 2791 37562
rect 2843 37510 2855 37562
rect 2907 37510 2919 37562
rect 2971 37510 6090 37562
rect 6142 37510 6154 37562
rect 6206 37510 6218 37562
rect 6270 37510 6282 37562
rect 6334 37510 6346 37562
rect 6398 37510 9517 37562
rect 9569 37510 9581 37562
rect 9633 37510 9645 37562
rect 9697 37510 9709 37562
rect 9761 37510 9773 37562
rect 9825 37510 12944 37562
rect 12996 37510 13008 37562
rect 13060 37510 13072 37562
rect 13124 37510 13136 37562
rect 13188 37510 13200 37562
rect 13252 37510 14812 37562
rect 1104 37488 14812 37510
rect 10778 37408 10784 37460
rect 10836 37408 10842 37460
rect 12618 37408 12624 37460
rect 12676 37408 12682 37460
rect 13173 37451 13231 37457
rect 13173 37417 13185 37451
rect 13219 37448 13231 37451
rect 13538 37448 13544 37460
rect 13219 37420 13544 37448
rect 13219 37417 13231 37420
rect 13173 37411 13231 37417
rect 13538 37408 13544 37420
rect 13596 37408 13602 37460
rect 12897 37383 12955 37389
rect 12897 37349 12909 37383
rect 12943 37349 12955 37383
rect 12897 37343 12955 37349
rect 1765 37315 1823 37321
rect 1765 37281 1777 37315
rect 1811 37312 1823 37315
rect 10502 37312 10508 37324
rect 1811 37284 10508 37312
rect 1811 37281 1823 37284
rect 1765 37275 1823 37281
rect 10502 37272 10508 37284
rect 10560 37312 10566 37324
rect 10560 37284 11008 37312
rect 10560 37272 10566 37284
rect 10980 37253 11008 37284
rect 10965 37247 11023 37253
rect 10965 37213 10977 37247
rect 11011 37213 11023 37247
rect 10965 37207 11023 37213
rect 12526 37204 12532 37256
rect 12584 37204 12590 37256
rect 12805 37247 12863 37253
rect 12805 37213 12817 37247
rect 12851 37244 12863 37247
rect 12912 37244 12940 37343
rect 13817 37315 13875 37321
rect 13817 37281 13829 37315
rect 13863 37312 13875 37315
rect 15378 37312 15384 37324
rect 13863 37284 15384 37312
rect 13863 37281 13875 37284
rect 13817 37275 13875 37281
rect 15378 37272 15384 37284
rect 15436 37272 15442 37324
rect 12851 37216 12940 37244
rect 12851 37213 12863 37216
rect 12805 37207 12863 37213
rect 13078 37204 13084 37256
rect 13136 37204 13142 37256
rect 13354 37204 13360 37256
rect 13412 37204 13418 37256
rect 14185 37247 14243 37253
rect 14185 37244 14197 37247
rect 13464 37216 14197 37244
rect 750 37136 756 37188
rect 808 37176 814 37188
rect 1489 37179 1547 37185
rect 1489 37176 1501 37179
rect 808 37148 1501 37176
rect 808 37136 814 37148
rect 1489 37145 1501 37148
rect 1535 37145 1547 37179
rect 1489 37139 1547 37145
rect 9122 37136 9128 37188
rect 9180 37176 9186 37188
rect 13464 37176 13492 37216
rect 14185 37213 14197 37216
rect 14231 37213 14243 37247
rect 14185 37207 14243 37213
rect 9180 37148 13492 37176
rect 13541 37179 13599 37185
rect 9180 37136 9186 37148
rect 13541 37145 13553 37179
rect 13587 37145 13599 37179
rect 13541 37139 13599 37145
rect 12342 37068 12348 37120
rect 12400 37068 12406 37120
rect 13078 37068 13084 37120
rect 13136 37108 13142 37120
rect 13556 37108 13584 37139
rect 13136 37080 13584 37108
rect 13136 37068 13142 37080
rect 14366 37068 14372 37120
rect 14424 37068 14430 37120
rect 1104 37018 14971 37040
rect 1104 36966 4376 37018
rect 4428 36966 4440 37018
rect 4492 36966 4504 37018
rect 4556 36966 4568 37018
rect 4620 36966 4632 37018
rect 4684 36966 7803 37018
rect 7855 36966 7867 37018
rect 7919 36966 7931 37018
rect 7983 36966 7995 37018
rect 8047 36966 8059 37018
rect 8111 36966 11230 37018
rect 11282 36966 11294 37018
rect 11346 36966 11358 37018
rect 11410 36966 11422 37018
rect 11474 36966 11486 37018
rect 11538 36966 14657 37018
rect 14709 36966 14721 37018
rect 14773 36966 14785 37018
rect 14837 36966 14849 37018
rect 14901 36966 14913 37018
rect 14965 36966 14971 37018
rect 1104 36944 14971 36966
rect 11885 36907 11943 36913
rect 11885 36873 11897 36907
rect 11931 36873 11943 36907
rect 12618 36904 12624 36916
rect 11885 36867 11943 36873
rect 12452 36876 12624 36904
rect 11900 36836 11928 36867
rect 12452 36836 12480 36876
rect 12618 36864 12624 36876
rect 12676 36864 12682 36916
rect 12713 36907 12771 36913
rect 12713 36873 12725 36907
rect 12759 36904 12771 36907
rect 13078 36904 13084 36916
rect 12759 36876 13084 36904
rect 12759 36873 12771 36876
rect 12713 36867 12771 36873
rect 13078 36864 13084 36876
rect 13136 36864 13142 36916
rect 14369 36907 14427 36913
rect 14369 36873 14381 36907
rect 14415 36873 14427 36907
rect 14369 36867 14427 36873
rect 11900 36808 12480 36836
rect 12544 36808 13216 36836
rect 11054 36728 11060 36780
rect 11112 36768 11118 36780
rect 12069 36771 12127 36777
rect 12069 36768 12081 36771
rect 11112 36740 12081 36768
rect 11112 36728 11118 36740
rect 12069 36737 12081 36740
rect 12115 36737 12127 36771
rect 12069 36731 12127 36737
rect 12158 36728 12164 36780
rect 12216 36768 12222 36780
rect 12345 36771 12403 36777
rect 12345 36768 12357 36771
rect 12216 36740 12357 36768
rect 12216 36728 12222 36740
rect 12345 36737 12357 36740
rect 12391 36737 12403 36771
rect 12544 36768 12572 36808
rect 12345 36731 12403 36737
rect 12452 36740 12572 36768
rect 12621 36771 12679 36777
rect 10134 36660 10140 36712
rect 10192 36700 10198 36712
rect 12452 36700 12480 36740
rect 12621 36737 12633 36771
rect 12667 36737 12679 36771
rect 12621 36731 12679 36737
rect 12636 36700 12664 36731
rect 12710 36728 12716 36780
rect 12768 36768 12774 36780
rect 13188 36777 13216 36808
rect 13630 36796 13636 36848
rect 13688 36836 13694 36848
rect 14384 36836 14412 36867
rect 13688 36808 14412 36836
rect 13688 36796 13694 36808
rect 12897 36771 12955 36777
rect 12897 36768 12909 36771
rect 12768 36740 12909 36768
rect 12768 36728 12774 36740
rect 12897 36737 12909 36740
rect 12943 36737 12955 36771
rect 12897 36731 12955 36737
rect 13173 36771 13231 36777
rect 13173 36737 13185 36771
rect 13219 36737 13231 36771
rect 13173 36731 13231 36737
rect 13541 36771 13599 36777
rect 13541 36737 13553 36771
rect 13587 36768 13599 36771
rect 13814 36768 13820 36780
rect 13587 36740 13820 36768
rect 13587 36737 13599 36740
rect 13541 36731 13599 36737
rect 13814 36728 13820 36740
rect 13872 36728 13878 36780
rect 13909 36771 13967 36777
rect 13909 36737 13921 36771
rect 13955 36768 13967 36771
rect 13998 36768 14004 36780
rect 13955 36740 14004 36768
rect 13955 36737 13967 36740
rect 13909 36731 13967 36737
rect 13998 36728 14004 36740
rect 14056 36728 14062 36780
rect 14093 36771 14151 36777
rect 14093 36737 14105 36771
rect 14139 36737 14151 36771
rect 14093 36731 14151 36737
rect 10192 36672 12480 36700
rect 12544 36672 12664 36700
rect 10192 36660 10198 36672
rect 12161 36635 12219 36641
rect 12161 36601 12173 36635
rect 12207 36632 12219 36635
rect 12250 36632 12256 36644
rect 12207 36604 12256 36632
rect 12207 36601 12219 36604
rect 12161 36595 12219 36601
rect 12250 36592 12256 36604
rect 12308 36592 12314 36644
rect 12342 36592 12348 36644
rect 12400 36632 12406 36644
rect 12544 36632 12572 36672
rect 13262 36660 13268 36712
rect 13320 36700 13326 36712
rect 14108 36700 14136 36731
rect 13320 36672 14136 36700
rect 13320 36660 13326 36672
rect 12400 36604 12572 36632
rect 12400 36592 12406 36604
rect 12434 36524 12440 36576
rect 12492 36524 12498 36576
rect 13722 36524 13728 36576
rect 13780 36524 13786 36576
rect 1104 36474 14812 36496
rect 1104 36422 2663 36474
rect 2715 36422 2727 36474
rect 2779 36422 2791 36474
rect 2843 36422 2855 36474
rect 2907 36422 2919 36474
rect 2971 36422 6090 36474
rect 6142 36422 6154 36474
rect 6206 36422 6218 36474
rect 6270 36422 6282 36474
rect 6334 36422 6346 36474
rect 6398 36422 9517 36474
rect 9569 36422 9581 36474
rect 9633 36422 9645 36474
rect 9697 36422 9709 36474
rect 9761 36422 9773 36474
rect 9825 36422 12944 36474
rect 12996 36422 13008 36474
rect 13060 36422 13072 36474
rect 13124 36422 13136 36474
rect 13188 36422 13200 36474
rect 13252 36422 14812 36474
rect 1104 36400 14812 36422
rect 9122 36320 9128 36372
rect 9180 36320 9186 36372
rect 11517 36363 11575 36369
rect 11517 36329 11529 36363
rect 11563 36360 11575 36363
rect 12158 36360 12164 36372
rect 11563 36332 12164 36360
rect 11563 36329 11575 36332
rect 11517 36323 11575 36329
rect 12158 36320 12164 36332
rect 12216 36320 12222 36372
rect 12342 36320 12348 36372
rect 12400 36320 12406 36372
rect 12621 36363 12679 36369
rect 12621 36329 12633 36363
rect 12667 36360 12679 36363
rect 12710 36360 12716 36372
rect 12667 36332 12716 36360
rect 12667 36329 12679 36332
rect 12621 36323 12679 36329
rect 12710 36320 12716 36332
rect 12768 36320 12774 36372
rect 13354 36320 13360 36372
rect 13412 36320 13418 36372
rect 11793 36295 11851 36301
rect 11793 36261 11805 36295
rect 11839 36292 11851 36295
rect 13372 36292 13400 36320
rect 11839 36264 13400 36292
rect 11839 36261 11851 36264
rect 11793 36255 11851 36261
rect 11808 36196 12848 36224
rect 11808 36168 11836 36196
rect 9306 36116 9312 36168
rect 9364 36116 9370 36168
rect 11701 36159 11759 36165
rect 11701 36156 11713 36159
rect 9416 36128 11713 36156
rect 750 36048 756 36100
rect 808 36088 814 36100
rect 1489 36091 1547 36097
rect 1489 36088 1501 36091
rect 808 36060 1501 36088
rect 808 36048 814 36060
rect 1489 36057 1501 36060
rect 1535 36057 1547 36091
rect 1489 36051 1547 36057
rect 1857 36091 1915 36097
rect 1857 36057 1869 36091
rect 1903 36088 1915 36091
rect 5810 36088 5816 36100
rect 1903 36060 5816 36088
rect 1903 36057 1915 36060
rect 1857 36051 1915 36057
rect 5810 36048 5816 36060
rect 5868 36088 5874 36100
rect 6822 36088 6828 36100
rect 5868 36060 6828 36088
rect 5868 36048 5874 36060
rect 6822 36048 6828 36060
rect 6880 36048 6886 36100
rect 8294 36048 8300 36100
rect 8352 36088 8358 36100
rect 9416 36088 9444 36128
rect 11701 36125 11713 36128
rect 11747 36125 11759 36159
rect 11701 36119 11759 36125
rect 11790 36116 11796 36168
rect 11848 36116 11854 36168
rect 11977 36159 12035 36165
rect 11977 36125 11989 36159
rect 12023 36125 12035 36159
rect 11977 36119 12035 36125
rect 8352 36060 9444 36088
rect 8352 36048 8358 36060
rect 7190 35980 7196 36032
rect 7248 36020 7254 36032
rect 11992 36020 12020 36119
rect 12158 36116 12164 36168
rect 12216 36156 12222 36168
rect 12820 36165 12848 36196
rect 12253 36159 12311 36165
rect 12253 36156 12265 36159
rect 12216 36128 12265 36156
rect 12216 36116 12222 36128
rect 12253 36125 12265 36128
rect 12299 36125 12311 36159
rect 12253 36119 12311 36125
rect 12529 36159 12587 36165
rect 12529 36125 12541 36159
rect 12575 36156 12587 36159
rect 12805 36159 12863 36165
rect 12575 36128 12756 36156
rect 12575 36125 12587 36128
rect 12529 36119 12587 36125
rect 12728 36100 12756 36128
rect 12805 36125 12817 36159
rect 12851 36125 12863 36159
rect 12805 36119 12863 36125
rect 14182 36116 14188 36168
rect 14240 36116 14246 36168
rect 12710 36048 12716 36100
rect 12768 36048 12774 36100
rect 12986 36048 12992 36100
rect 13044 36048 13050 36100
rect 13170 36048 13176 36100
rect 13228 36088 13234 36100
rect 13541 36091 13599 36097
rect 13541 36088 13553 36091
rect 13228 36060 13553 36088
rect 13228 36048 13234 36060
rect 13541 36057 13553 36060
rect 13587 36057 13599 36091
rect 13541 36051 13599 36057
rect 13909 36091 13967 36097
rect 13909 36057 13921 36091
rect 13955 36088 13967 36091
rect 15562 36088 15568 36100
rect 13955 36060 15568 36088
rect 13955 36057 13967 36060
rect 13909 36051 13967 36057
rect 15562 36048 15568 36060
rect 15620 36048 15626 36100
rect 7248 35992 12020 36020
rect 7248 35980 7254 35992
rect 12066 35980 12072 36032
rect 12124 35980 12130 36032
rect 13262 35980 13268 36032
rect 13320 35980 13326 36032
rect 14369 36023 14427 36029
rect 14369 35989 14381 36023
rect 14415 36020 14427 36023
rect 15102 36020 15108 36032
rect 14415 35992 15108 36020
rect 14415 35989 14427 35992
rect 14369 35983 14427 35989
rect 15102 35980 15108 35992
rect 15160 35980 15166 36032
rect 1104 35930 14971 35952
rect 1104 35878 4376 35930
rect 4428 35878 4440 35930
rect 4492 35878 4504 35930
rect 4556 35878 4568 35930
rect 4620 35878 4632 35930
rect 4684 35878 7803 35930
rect 7855 35878 7867 35930
rect 7919 35878 7931 35930
rect 7983 35878 7995 35930
rect 8047 35878 8059 35930
rect 8111 35878 11230 35930
rect 11282 35878 11294 35930
rect 11346 35878 11358 35930
rect 11410 35878 11422 35930
rect 11474 35878 11486 35930
rect 11538 35878 14657 35930
rect 14709 35878 14721 35930
rect 14773 35878 14785 35930
rect 14837 35878 14849 35930
rect 14901 35878 14913 35930
rect 14965 35878 14971 35930
rect 1104 35856 14971 35878
rect 1762 35776 1768 35828
rect 1820 35776 1826 35828
rect 8389 35819 8447 35825
rect 8389 35785 8401 35819
rect 8435 35816 8447 35819
rect 9306 35816 9312 35828
rect 8435 35788 9312 35816
rect 8435 35785 8447 35788
rect 8389 35779 8447 35785
rect 9306 35776 9312 35788
rect 9364 35776 9370 35828
rect 10134 35776 10140 35828
rect 10192 35776 10198 35828
rect 11517 35819 11575 35825
rect 11517 35785 11529 35819
rect 11563 35785 11575 35819
rect 11517 35779 11575 35785
rect 11793 35819 11851 35825
rect 11793 35785 11805 35819
rect 11839 35816 11851 35819
rect 11839 35788 13032 35816
rect 11839 35785 11851 35788
rect 11793 35779 11851 35785
rect 10226 35708 10232 35760
rect 10284 35748 10290 35760
rect 11532 35748 11560 35779
rect 10284 35720 11468 35748
rect 11532 35720 12388 35748
rect 10284 35708 10290 35720
rect 750 35640 756 35692
rect 808 35680 814 35692
rect 1397 35683 1455 35689
rect 1397 35680 1409 35683
rect 808 35652 1409 35680
rect 808 35640 814 35652
rect 1397 35649 1409 35652
rect 1443 35649 1455 35683
rect 1397 35643 1455 35649
rect 1946 35640 1952 35692
rect 2004 35640 2010 35692
rect 8570 35640 8576 35692
rect 8628 35640 8634 35692
rect 10318 35640 10324 35692
rect 10376 35640 10382 35692
rect 11333 35683 11391 35689
rect 11333 35649 11345 35683
rect 11379 35649 11391 35683
rect 11333 35643 11391 35649
rect 11149 35547 11207 35553
rect 11149 35513 11161 35547
rect 11195 35513 11207 35547
rect 11348 35544 11376 35643
rect 11440 35612 11468 35720
rect 11701 35683 11759 35689
rect 11701 35649 11713 35683
rect 11747 35680 11759 35683
rect 11882 35680 11888 35692
rect 11747 35652 11888 35680
rect 11747 35649 11759 35652
rect 11701 35643 11759 35649
rect 11882 35640 11888 35652
rect 11940 35640 11946 35692
rect 11977 35683 12035 35689
rect 11977 35649 11989 35683
rect 12023 35649 12035 35683
rect 11977 35643 12035 35649
rect 11992 35612 12020 35643
rect 12066 35640 12072 35692
rect 12124 35684 12130 35692
rect 12124 35680 12202 35684
rect 12253 35683 12311 35689
rect 12253 35680 12265 35683
rect 12124 35656 12265 35680
rect 12124 35640 12130 35656
rect 12174 35652 12265 35656
rect 12253 35649 12265 35652
rect 12299 35649 12311 35683
rect 12360 35680 12388 35720
rect 12434 35708 12440 35760
rect 12492 35708 12498 35760
rect 13004 35757 13032 35788
rect 14182 35776 14188 35828
rect 14240 35776 14246 35828
rect 12989 35751 13047 35757
rect 12989 35717 13001 35751
rect 13035 35717 13047 35751
rect 14200 35748 14228 35776
rect 12989 35711 13047 35717
rect 13096 35720 14228 35748
rect 13096 35680 13124 35720
rect 12360 35652 13124 35680
rect 13357 35683 13415 35689
rect 12253 35643 12311 35649
rect 13357 35649 13369 35683
rect 13403 35649 13415 35683
rect 13357 35643 13415 35649
rect 13170 35612 13176 35624
rect 11440 35584 12020 35612
rect 12406 35584 13176 35612
rect 12069 35547 12127 35553
rect 12069 35544 12081 35547
rect 11348 35516 12081 35544
rect 11149 35507 11207 35513
rect 12069 35513 12081 35516
rect 12115 35513 12127 35547
rect 12069 35507 12127 35513
rect 1581 35479 1639 35485
rect 1581 35445 1593 35479
rect 1627 35476 1639 35479
rect 5994 35476 6000 35488
rect 1627 35448 6000 35476
rect 1627 35445 1639 35448
rect 1581 35439 1639 35445
rect 5994 35436 6000 35448
rect 6052 35436 6058 35488
rect 11164 35476 11192 35507
rect 12406 35476 12434 35584
rect 13170 35572 13176 35584
rect 13228 35572 13234 35624
rect 13372 35612 13400 35643
rect 13538 35640 13544 35692
rect 13596 35640 13602 35692
rect 13630 35640 13636 35692
rect 13688 35680 13694 35692
rect 14093 35683 14151 35689
rect 14093 35680 14105 35683
rect 13688 35652 14105 35680
rect 13688 35640 13694 35652
rect 14093 35649 14105 35652
rect 14139 35649 14151 35683
rect 14093 35643 14151 35649
rect 14458 35612 14464 35624
rect 13372 35584 14464 35612
rect 14458 35572 14464 35584
rect 14516 35572 14522 35624
rect 15102 35544 15108 35556
rect 12728 35516 15108 35544
rect 12728 35485 12756 35516
rect 15102 35504 15108 35516
rect 15160 35504 15166 35556
rect 11164 35448 12434 35476
rect 12713 35479 12771 35485
rect 12713 35445 12725 35479
rect 12759 35445 12771 35479
rect 12713 35439 12771 35445
rect 13814 35436 13820 35488
rect 13872 35436 13878 35488
rect 14369 35479 14427 35485
rect 14369 35445 14381 35479
rect 14415 35476 14427 35479
rect 15470 35476 15476 35488
rect 14415 35448 15476 35476
rect 14415 35445 14427 35448
rect 14369 35439 14427 35445
rect 15470 35436 15476 35448
rect 15528 35436 15534 35488
rect 1104 35386 14812 35408
rect 1104 35334 2663 35386
rect 2715 35334 2727 35386
rect 2779 35334 2791 35386
rect 2843 35334 2855 35386
rect 2907 35334 2919 35386
rect 2971 35334 6090 35386
rect 6142 35334 6154 35386
rect 6206 35334 6218 35386
rect 6270 35334 6282 35386
rect 6334 35334 6346 35386
rect 6398 35334 9517 35386
rect 9569 35334 9581 35386
rect 9633 35334 9645 35386
rect 9697 35334 9709 35386
rect 9761 35334 9773 35386
rect 9825 35334 12944 35386
rect 12996 35334 13008 35386
rect 13060 35334 13072 35386
rect 13124 35334 13136 35386
rect 13188 35334 13200 35386
rect 13252 35334 14812 35386
rect 1104 35312 14812 35334
rect 1581 35275 1639 35281
rect 1581 35241 1593 35275
rect 1627 35272 1639 35275
rect 1946 35272 1952 35284
rect 1627 35244 1952 35272
rect 1627 35241 1639 35244
rect 1581 35235 1639 35241
rect 1946 35232 1952 35244
rect 2004 35232 2010 35284
rect 9309 35275 9367 35281
rect 9309 35241 9321 35275
rect 9355 35272 9367 35275
rect 10318 35272 10324 35284
rect 9355 35244 10324 35272
rect 9355 35241 9367 35244
rect 9309 35235 9367 35241
rect 10318 35232 10324 35244
rect 10376 35232 10382 35284
rect 11241 35275 11299 35281
rect 11241 35241 11253 35275
rect 11287 35272 11299 35275
rect 12802 35272 12808 35284
rect 11287 35244 12808 35272
rect 11287 35241 11299 35244
rect 11241 35235 11299 35241
rect 12802 35232 12808 35244
rect 12860 35232 12866 35284
rect 12912 35244 14320 35272
rect 6822 35096 6828 35148
rect 6880 35136 6886 35148
rect 11054 35136 11060 35148
rect 6880 35108 11060 35136
rect 6880 35096 6886 35108
rect 11054 35096 11060 35108
rect 11112 35096 11118 35148
rect 11514 35096 11520 35148
rect 11572 35096 11578 35148
rect 1765 35071 1823 35077
rect 1765 35037 1777 35071
rect 1811 35037 1823 35071
rect 1765 35031 1823 35037
rect 1780 35000 1808 35031
rect 5534 35028 5540 35080
rect 5592 35068 5598 35080
rect 9493 35071 9551 35077
rect 9493 35068 9505 35071
rect 5592 35040 9505 35068
rect 5592 35028 5598 35040
rect 9493 35037 9505 35040
rect 9539 35037 9551 35071
rect 9493 35031 9551 35037
rect 10962 35028 10968 35080
rect 11020 35068 11026 35080
rect 11425 35071 11483 35077
rect 11425 35068 11437 35071
rect 11020 35040 11437 35068
rect 11020 35028 11026 35040
rect 11425 35037 11437 35040
rect 11471 35037 11483 35071
rect 11759 35071 11817 35077
rect 11759 35068 11771 35071
rect 11425 35031 11483 35037
rect 11532 35040 11771 35068
rect 6914 35000 6920 35012
rect 1780 34972 6920 35000
rect 6914 34960 6920 34972
rect 6972 34960 6978 35012
rect 11146 34960 11152 35012
rect 11204 35000 11210 35012
rect 11532 35000 11560 35040
rect 11759 35037 11771 35040
rect 11805 35068 11817 35071
rect 12158 35068 12164 35080
rect 11805 35040 12164 35068
rect 11805 35037 11817 35040
rect 11759 35031 11817 35037
rect 12158 35028 12164 35040
rect 12216 35028 12222 35080
rect 12912 35068 12940 35244
rect 14093 35207 14151 35213
rect 14093 35173 14105 35207
rect 14139 35173 14151 35207
rect 14093 35167 14151 35173
rect 12268 35040 12940 35068
rect 12989 35071 13047 35077
rect 11204 34972 11560 35000
rect 11204 34960 11210 34972
rect 10410 34892 10416 34944
rect 10468 34932 10474 34944
rect 12268 34932 12296 35040
rect 12989 35037 13001 35071
rect 13035 35064 13047 35071
rect 14108 35068 14136 35167
rect 14292 35077 14320 35244
rect 13096 35064 14136 35068
rect 13035 35040 14136 35064
rect 14277 35071 14335 35077
rect 13035 35037 13124 35040
rect 12989 35036 13124 35037
rect 14277 35037 14289 35071
rect 14323 35037 14335 35071
rect 12989 35031 13047 35036
rect 14277 35031 14335 35037
rect 13541 35003 13599 35009
rect 13541 35000 13553 35003
rect 12406 34972 13553 35000
rect 12406 34944 12434 34972
rect 13541 34969 13553 34972
rect 13587 34969 13599 35003
rect 13541 34963 13599 34969
rect 13909 35003 13967 35009
rect 13909 34969 13921 35003
rect 13955 35000 13967 35003
rect 14550 35000 14556 35012
rect 13955 34972 14556 35000
rect 13955 34969 13967 34972
rect 13909 34963 13967 34969
rect 14550 34960 14556 34972
rect 14608 34960 14614 35012
rect 10468 34904 12296 34932
rect 10468 34892 10474 34904
rect 12342 34892 12348 34944
rect 12400 34904 12434 34944
rect 12400 34892 12406 34904
rect 12526 34892 12532 34944
rect 12584 34892 12590 34944
rect 13262 34892 13268 34944
rect 13320 34892 13326 34944
rect 1104 34842 14971 34864
rect 1104 34790 4376 34842
rect 4428 34790 4440 34842
rect 4492 34790 4504 34842
rect 4556 34790 4568 34842
rect 4620 34790 4632 34842
rect 4684 34790 7803 34842
rect 7855 34790 7867 34842
rect 7919 34790 7931 34842
rect 7983 34790 7995 34842
rect 8047 34790 8059 34842
rect 8111 34790 11230 34842
rect 11282 34790 11294 34842
rect 11346 34790 11358 34842
rect 11410 34790 11422 34842
rect 11474 34790 11486 34842
rect 11538 34790 14657 34842
rect 14709 34790 14721 34842
rect 14773 34790 14785 34842
rect 14837 34790 14849 34842
rect 14901 34790 14913 34842
rect 14965 34790 14971 34842
rect 1104 34768 14971 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 5718 34728 5724 34740
rect 1627 34700 5724 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 5718 34688 5724 34700
rect 5776 34728 5782 34740
rect 6822 34728 6828 34740
rect 5776 34700 6828 34728
rect 5776 34688 5782 34700
rect 6822 34688 6828 34700
rect 6880 34688 6886 34740
rect 10410 34688 10416 34740
rect 10468 34688 10474 34740
rect 10689 34731 10747 34737
rect 10689 34697 10701 34731
rect 10735 34697 10747 34731
rect 10689 34691 10747 34697
rect 10704 34660 10732 34691
rect 10962 34688 10968 34740
rect 11020 34688 11026 34740
rect 11517 34731 11575 34737
rect 11517 34697 11529 34731
rect 11563 34728 11575 34731
rect 13538 34728 13544 34740
rect 11563 34700 13544 34728
rect 11563 34697 11575 34700
rect 11517 34691 11575 34697
rect 13538 34688 13544 34700
rect 13596 34688 13602 34740
rect 11885 34663 11943 34669
rect 11885 34660 11897 34663
rect 10704 34632 11897 34660
rect 11885 34629 11897 34632
rect 11931 34629 11943 34663
rect 11885 34623 11943 34629
rect 11974 34620 11980 34672
rect 12032 34660 12038 34672
rect 12989 34663 13047 34669
rect 12989 34660 13001 34663
rect 12032 34632 13001 34660
rect 12032 34620 12038 34632
rect 12989 34629 13001 34632
rect 13035 34629 13047 34663
rect 12989 34623 13047 34629
rect 1394 34552 1400 34604
rect 1452 34552 1458 34604
rect 10594 34552 10600 34604
rect 10652 34552 10658 34604
rect 10870 34552 10876 34604
rect 10928 34552 10934 34604
rect 11054 34552 11060 34604
rect 11112 34592 11118 34604
rect 11149 34595 11207 34601
rect 11149 34592 11161 34595
rect 11112 34564 11161 34592
rect 11112 34552 11118 34564
rect 11149 34561 11161 34564
rect 11195 34561 11207 34595
rect 11149 34555 11207 34561
rect 11701 34595 11759 34601
rect 11701 34561 11713 34595
rect 11747 34561 11759 34595
rect 11701 34555 11759 34561
rect 10502 34484 10508 34536
rect 10560 34524 10566 34536
rect 11716 34524 11744 34555
rect 12250 34552 12256 34604
rect 12308 34552 12314 34604
rect 12434 34552 12440 34604
rect 12492 34552 12498 34604
rect 13354 34552 13360 34604
rect 13412 34552 13418 34604
rect 13538 34552 13544 34604
rect 13596 34552 13602 34604
rect 14090 34552 14096 34604
rect 14148 34552 14154 34604
rect 14461 34595 14519 34601
rect 14461 34561 14473 34595
rect 14507 34592 14519 34595
rect 15654 34592 15660 34604
rect 14507 34564 15660 34592
rect 14507 34561 14519 34564
rect 14461 34555 14519 34561
rect 15654 34552 15660 34564
rect 15712 34552 15718 34604
rect 10560 34496 11744 34524
rect 10560 34484 10566 34496
rect 12342 34484 12348 34536
rect 12400 34524 12406 34536
rect 12713 34527 12771 34533
rect 12713 34524 12725 34527
rect 12400 34496 12725 34524
rect 12400 34484 12406 34496
rect 12713 34493 12725 34496
rect 12759 34493 12771 34527
rect 12713 34487 12771 34493
rect 13814 34348 13820 34400
rect 13872 34348 13878 34400
rect 1104 34298 14812 34320
rect 1104 34246 2663 34298
rect 2715 34246 2727 34298
rect 2779 34246 2791 34298
rect 2843 34246 2855 34298
rect 2907 34246 2919 34298
rect 2971 34246 6090 34298
rect 6142 34246 6154 34298
rect 6206 34246 6218 34298
rect 6270 34246 6282 34298
rect 6334 34246 6346 34298
rect 6398 34246 9517 34298
rect 9569 34246 9581 34298
rect 9633 34246 9645 34298
rect 9697 34246 9709 34298
rect 9761 34246 9773 34298
rect 9825 34246 12944 34298
rect 12996 34246 13008 34298
rect 13060 34246 13072 34298
rect 13124 34246 13136 34298
rect 13188 34246 13200 34298
rect 13252 34246 14812 34298
rect 1104 34224 14812 34246
rect 10226 34144 10232 34196
rect 10284 34144 10290 34196
rect 10502 34144 10508 34196
rect 10560 34144 10566 34196
rect 11606 34008 11612 34060
rect 11664 34048 11670 34060
rect 12161 34051 12219 34057
rect 12161 34048 12173 34051
rect 11664 34020 12173 34048
rect 11664 34008 11670 34020
rect 12161 34017 12173 34020
rect 12207 34017 12219 34051
rect 12161 34011 12219 34017
rect 750 33940 756 33992
rect 808 33980 814 33992
rect 1397 33983 1455 33989
rect 1397 33980 1409 33983
rect 808 33952 1409 33980
rect 808 33940 814 33952
rect 1397 33949 1409 33952
rect 1443 33949 1455 33983
rect 1397 33943 1455 33949
rect 8754 33940 8760 33992
rect 8812 33980 8818 33992
rect 10413 33983 10471 33989
rect 10413 33980 10425 33983
rect 8812 33952 10425 33980
rect 8812 33940 8818 33952
rect 10413 33949 10425 33952
rect 10459 33949 10471 33983
rect 10413 33943 10471 33949
rect 10689 33983 10747 33989
rect 10689 33949 10701 33983
rect 10735 33949 10747 33983
rect 10689 33943 10747 33949
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33949 10839 33983
rect 10781 33943 10839 33949
rect 11055 33983 11113 33989
rect 11055 33949 11067 33983
rect 11101 33980 11113 33983
rect 11514 33980 11520 33992
rect 11101 33952 11520 33980
rect 11101 33949 11113 33952
rect 11055 33943 11113 33949
rect 10704 33912 10732 33943
rect 10336 33884 10732 33912
rect 10796 33912 10824 33943
rect 11514 33940 11520 33952
rect 11572 33980 11578 33992
rect 11790 33980 11796 33992
rect 11572 33952 11796 33980
rect 11572 33940 11578 33952
rect 11790 33940 11796 33952
rect 11848 33940 11854 33992
rect 12802 33980 12808 33992
rect 12418 33979 12808 33980
rect 12403 33973 12808 33979
rect 12403 33970 12415 33973
rect 12314 33942 12415 33970
rect 11606 33912 11612 33924
rect 10796 33884 11612 33912
rect 10336 33856 10364 33884
rect 11606 33872 11612 33884
rect 11664 33872 11670 33924
rect 12314 33912 12342 33942
rect 12403 33939 12415 33942
rect 12449 33952 12808 33973
rect 12449 33939 12461 33952
rect 12802 33940 12808 33952
rect 12860 33940 12866 33992
rect 12986 33940 12992 33992
rect 13044 33980 13050 33992
rect 13725 33983 13783 33989
rect 13725 33980 13737 33983
rect 13044 33952 13737 33980
rect 13044 33940 13050 33952
rect 13725 33949 13737 33952
rect 13771 33949 13783 33983
rect 13725 33943 13783 33949
rect 14274 33940 14280 33992
rect 14332 33940 14338 33992
rect 12403 33933 12461 33939
rect 11716 33884 12342 33912
rect 1581 33847 1639 33853
rect 1581 33813 1593 33847
rect 1627 33844 1639 33847
rect 3602 33844 3608 33856
rect 1627 33816 3608 33844
rect 1627 33813 1639 33816
rect 1581 33807 1639 33813
rect 3602 33804 3608 33816
rect 3660 33844 3666 33856
rect 9858 33844 9864 33856
rect 3660 33816 9864 33844
rect 3660 33804 3666 33816
rect 9858 33804 9864 33816
rect 9916 33804 9922 33856
rect 10318 33804 10324 33856
rect 10376 33804 10382 33856
rect 10502 33804 10508 33856
rect 10560 33844 10566 33856
rect 11716 33844 11744 33884
rect 12710 33872 12716 33924
rect 12768 33912 12774 33924
rect 12768 33884 14136 33912
rect 12768 33872 12774 33884
rect 10560 33816 11744 33844
rect 11793 33847 11851 33853
rect 10560 33804 10566 33816
rect 11793 33813 11805 33847
rect 11839 33844 11851 33847
rect 12066 33844 12072 33856
rect 11839 33816 12072 33844
rect 11839 33813 11851 33816
rect 11793 33807 11851 33813
rect 12066 33804 12072 33816
rect 12124 33804 12130 33856
rect 13173 33847 13231 33853
rect 13173 33813 13185 33847
rect 13219 33844 13231 33847
rect 13262 33844 13268 33856
rect 13219 33816 13268 33844
rect 13219 33813 13231 33816
rect 13173 33807 13231 33813
rect 13262 33804 13268 33816
rect 13320 33804 13326 33856
rect 13538 33804 13544 33856
rect 13596 33804 13602 33856
rect 14108 33853 14136 33884
rect 14093 33847 14151 33853
rect 14093 33813 14105 33847
rect 14139 33813 14151 33847
rect 14093 33807 14151 33813
rect 1104 33754 14971 33776
rect 1104 33702 4376 33754
rect 4428 33702 4440 33754
rect 4492 33702 4504 33754
rect 4556 33702 4568 33754
rect 4620 33702 4632 33754
rect 4684 33702 7803 33754
rect 7855 33702 7867 33754
rect 7919 33702 7931 33754
rect 7983 33702 7995 33754
rect 8047 33702 8059 33754
rect 8111 33702 11230 33754
rect 11282 33702 11294 33754
rect 11346 33702 11358 33754
rect 11410 33702 11422 33754
rect 11474 33702 11486 33754
rect 11538 33702 14657 33754
rect 14709 33702 14721 33754
rect 14773 33702 14785 33754
rect 14837 33702 14849 33754
rect 14901 33702 14913 33754
rect 14965 33702 14971 33754
rect 1104 33680 14971 33702
rect 11609 33643 11667 33649
rect 11609 33609 11621 33643
rect 11655 33640 11667 33643
rect 12158 33640 12164 33652
rect 11655 33612 12164 33640
rect 11655 33609 11667 33612
rect 11609 33603 11667 33609
rect 12158 33600 12164 33612
rect 12216 33600 12222 33652
rect 10778 33532 10784 33584
rect 10836 33572 10842 33584
rect 13541 33575 13599 33581
rect 13541 33572 13553 33575
rect 10836 33544 13553 33572
rect 10836 33532 10842 33544
rect 13541 33541 13553 33544
rect 13587 33541 13599 33575
rect 13541 33535 13599 33541
rect 11790 33464 11796 33516
rect 11848 33464 11854 33516
rect 12158 33504 12164 33516
rect 12071 33476 12164 33504
rect 12158 33464 12164 33476
rect 12216 33504 12222 33516
rect 13998 33504 14004 33516
rect 12216 33476 14004 33504
rect 12216 33464 12222 33476
rect 13998 33464 14004 33476
rect 14056 33464 14062 33516
rect 14093 33507 14151 33513
rect 14093 33473 14105 33507
rect 14139 33504 14151 33507
rect 15378 33504 15384 33516
rect 14139 33476 15384 33504
rect 14139 33473 14151 33476
rect 14093 33467 14151 33473
rect 15378 33464 15384 33476
rect 15436 33464 15442 33516
rect 11606 33396 11612 33448
rect 11664 33436 11670 33448
rect 11885 33439 11943 33445
rect 11885 33436 11897 33439
rect 11664 33408 11897 33436
rect 11664 33396 11670 33408
rect 11885 33405 11897 33408
rect 11931 33405 11943 33439
rect 11885 33399 11943 33405
rect 12544 33340 13032 33368
rect 10134 33260 10140 33312
rect 10192 33300 10198 33312
rect 12544 33300 12572 33340
rect 13004 33312 13032 33340
rect 10192 33272 12572 33300
rect 10192 33260 10198 33272
rect 12894 33260 12900 33312
rect 12952 33260 12958 33312
rect 12986 33260 12992 33312
rect 13044 33260 13050 33312
rect 13817 33303 13875 33309
rect 13817 33269 13829 33303
rect 13863 33300 13875 33303
rect 13998 33300 14004 33312
rect 13863 33272 14004 33300
rect 13863 33269 13875 33272
rect 13817 33263 13875 33269
rect 13998 33260 14004 33272
rect 14056 33260 14062 33312
rect 14182 33260 14188 33312
rect 14240 33260 14246 33312
rect 1104 33210 14812 33232
rect 1104 33158 2663 33210
rect 2715 33158 2727 33210
rect 2779 33158 2791 33210
rect 2843 33158 2855 33210
rect 2907 33158 2919 33210
rect 2971 33158 6090 33210
rect 6142 33158 6154 33210
rect 6206 33158 6218 33210
rect 6270 33158 6282 33210
rect 6334 33158 6346 33210
rect 6398 33158 9517 33210
rect 9569 33158 9581 33210
rect 9633 33158 9645 33210
rect 9697 33158 9709 33210
rect 9761 33158 9773 33210
rect 9825 33158 12944 33210
rect 12996 33158 13008 33210
rect 13060 33158 13072 33210
rect 13124 33158 13136 33210
rect 13188 33158 13200 33210
rect 13252 33158 14812 33210
rect 1104 33136 14812 33158
rect 9493 33099 9551 33105
rect 9493 33065 9505 33099
rect 9539 33096 9551 33099
rect 10042 33096 10048 33108
rect 9539 33068 10048 33096
rect 9539 33065 9551 33068
rect 9493 33059 9551 33065
rect 10042 33056 10048 33068
rect 10100 33056 10106 33108
rect 10505 33099 10563 33105
rect 10505 33065 10517 33099
rect 10551 33096 10563 33099
rect 10686 33096 10692 33108
rect 10551 33068 10692 33096
rect 10551 33065 10563 33068
rect 10505 33059 10563 33065
rect 10686 33056 10692 33068
rect 10744 33056 10750 33108
rect 11241 33099 11299 33105
rect 11241 33065 11253 33099
rect 11287 33096 11299 33099
rect 11790 33096 11796 33108
rect 11287 33068 11796 33096
rect 11287 33065 11299 33068
rect 11241 33059 11299 33065
rect 11790 33056 11796 33068
rect 11848 33056 11854 33108
rect 12434 33056 12440 33108
rect 12492 33096 12498 33108
rect 14093 33099 14151 33105
rect 14093 33096 14105 33099
rect 12492 33068 14105 33096
rect 12492 33056 12498 33068
rect 14093 33065 14105 33068
rect 14139 33065 14151 33099
rect 14093 33059 14151 33065
rect 9953 33031 10011 33037
rect 9953 32997 9965 33031
rect 9999 32997 10011 33031
rect 9953 32991 10011 32997
rect 10965 33031 11023 33037
rect 10965 32997 10977 33031
rect 11011 33028 11023 33031
rect 11011 33000 12434 33028
rect 11011 32997 11023 33000
rect 10965 32991 11023 32997
rect 9968 32960 9996 32991
rect 9968 32932 10732 32960
rect 750 32852 756 32904
rect 808 32892 814 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 808 32864 1409 32892
rect 808 32852 814 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 8938 32852 8944 32904
rect 8996 32892 9002 32904
rect 10704 32901 10732 32932
rect 10870 32920 10876 32972
rect 10928 32920 10934 32972
rect 9677 32895 9735 32901
rect 9677 32892 9689 32895
rect 8996 32864 9689 32892
rect 8996 32852 9002 32864
rect 9677 32861 9689 32864
rect 9723 32861 9735 32895
rect 9677 32855 9735 32861
rect 10137 32895 10195 32901
rect 10137 32861 10149 32895
rect 10183 32861 10195 32895
rect 10137 32855 10195 32861
rect 10689 32895 10747 32901
rect 10689 32861 10701 32895
rect 10735 32861 10747 32895
rect 10689 32855 10747 32861
rect 8478 32784 8484 32836
rect 8536 32824 8542 32836
rect 10152 32824 10180 32855
rect 8536 32796 10180 32824
rect 8536 32784 8542 32796
rect 1581 32759 1639 32765
rect 1581 32725 1593 32759
rect 1627 32756 1639 32759
rect 6454 32756 6460 32768
rect 1627 32728 6460 32756
rect 1627 32725 1639 32728
rect 1581 32719 1639 32725
rect 6454 32716 6460 32728
rect 6512 32716 6518 32768
rect 7282 32716 7288 32768
rect 7340 32756 7346 32768
rect 10888 32756 10916 32920
rect 11146 32852 11152 32904
rect 11204 32852 11210 32904
rect 11425 32895 11483 32901
rect 11425 32861 11437 32895
rect 11471 32861 11483 32895
rect 11425 32855 11483 32861
rect 11701 32895 11759 32901
rect 11701 32861 11713 32895
rect 11747 32892 11759 32895
rect 12406 32892 12434 33000
rect 13722 32988 13728 33040
rect 13780 33028 13786 33040
rect 14274 33028 14280 33040
rect 13780 33000 14280 33028
rect 13780 32988 13786 33000
rect 14274 32988 14280 33000
rect 14332 32988 14338 33040
rect 12713 32963 12771 32969
rect 12713 32929 12725 32963
rect 12759 32960 12771 32963
rect 15562 32960 15568 32972
rect 12759 32932 15568 32960
rect 12759 32929 12771 32932
rect 12713 32923 12771 32929
rect 15562 32920 15568 32932
rect 15620 32920 15626 32972
rect 12989 32895 13047 32901
rect 12989 32892 13001 32895
rect 11747 32864 12342 32892
rect 12406 32864 13001 32892
rect 11747 32861 11759 32864
rect 11701 32855 11759 32861
rect 11440 32824 11468 32855
rect 11072 32796 11468 32824
rect 11072 32768 11100 32796
rect 11882 32784 11888 32836
rect 11940 32784 11946 32836
rect 7340 32728 10916 32756
rect 7340 32716 7346 32728
rect 11054 32716 11060 32768
rect 11112 32716 11118 32768
rect 11517 32759 11575 32765
rect 11517 32725 11529 32759
rect 11563 32756 11575 32759
rect 11974 32756 11980 32768
rect 11563 32728 11980 32756
rect 11563 32725 11575 32728
rect 11517 32719 11575 32725
rect 11974 32716 11980 32728
rect 12032 32716 12038 32768
rect 12158 32716 12164 32768
rect 12216 32716 12222 32768
rect 12314 32756 12342 32864
rect 12989 32861 13001 32864
rect 13035 32861 13047 32895
rect 12989 32855 13047 32861
rect 14274 32852 14280 32904
rect 14332 32852 14338 32904
rect 12434 32784 12440 32836
rect 12492 32784 12498 32836
rect 12710 32784 12716 32836
rect 12768 32784 12774 32836
rect 13354 32784 13360 32836
rect 13412 32784 13418 32836
rect 13541 32827 13599 32833
rect 13541 32793 13553 32827
rect 13587 32793 13599 32827
rect 13541 32787 13599 32793
rect 13909 32827 13967 32833
rect 13909 32793 13921 32827
rect 13955 32824 13967 32827
rect 14550 32824 14556 32836
rect 13955 32796 14556 32824
rect 13955 32793 13967 32796
rect 13909 32787 13967 32793
rect 12728 32756 12756 32784
rect 12314 32728 12756 32756
rect 12986 32716 12992 32768
rect 13044 32756 13050 32768
rect 13556 32756 13584 32787
rect 14550 32784 14556 32796
rect 14608 32784 14614 32836
rect 13044 32728 13584 32756
rect 13044 32716 13050 32728
rect 1104 32666 14971 32688
rect 1104 32614 4376 32666
rect 4428 32614 4440 32666
rect 4492 32614 4504 32666
rect 4556 32614 4568 32666
rect 4620 32614 4632 32666
rect 4684 32614 7803 32666
rect 7855 32614 7867 32666
rect 7919 32614 7931 32666
rect 7983 32614 7995 32666
rect 8047 32614 8059 32666
rect 8111 32614 11230 32666
rect 11282 32614 11294 32666
rect 11346 32614 11358 32666
rect 11410 32614 11422 32666
rect 11474 32614 11486 32666
rect 11538 32614 14657 32666
rect 14709 32614 14721 32666
rect 14773 32614 14785 32666
rect 14837 32614 14849 32666
rect 14901 32614 14913 32666
rect 14965 32614 14971 32666
rect 1104 32592 14971 32614
rect 2041 32555 2099 32561
rect 2041 32521 2053 32555
rect 2087 32552 2099 32555
rect 2222 32552 2228 32564
rect 2087 32524 2228 32552
rect 2087 32521 2099 32524
rect 2041 32515 2099 32521
rect 2222 32512 2228 32524
rect 2280 32512 2286 32564
rect 7024 32524 8432 32552
rect 750 32376 756 32428
rect 808 32416 814 32428
rect 1397 32419 1455 32425
rect 1397 32416 1409 32419
rect 808 32388 1409 32416
rect 808 32376 814 32388
rect 1397 32385 1409 32388
rect 1443 32385 1455 32419
rect 1397 32379 1455 32385
rect 2222 32376 2228 32428
rect 2280 32376 2286 32428
rect 6914 32376 6920 32428
rect 6972 32416 6978 32428
rect 7024 32425 7052 32524
rect 7267 32449 7325 32455
rect 7009 32419 7067 32425
rect 7009 32416 7021 32419
rect 6972 32388 7021 32416
rect 6972 32376 6978 32388
rect 7009 32385 7021 32388
rect 7055 32385 7067 32419
rect 7267 32415 7279 32449
rect 7313 32446 7325 32449
rect 7313 32428 7328 32446
rect 7267 32409 7288 32415
rect 7009 32379 7067 32385
rect 7282 32376 7288 32409
rect 7340 32376 7346 32428
rect 8404 32425 8432 32524
rect 8662 32512 8668 32564
rect 8720 32552 8726 32564
rect 8720 32524 9812 32552
rect 8720 32512 8726 32524
rect 8478 32444 8484 32496
rect 8536 32484 8542 32496
rect 8536 32456 8616 32484
rect 8536 32444 8542 32456
rect 8588 32446 8616 32456
rect 8647 32449 8705 32455
rect 8647 32446 8659 32449
rect 8389 32419 8447 32425
rect 8389 32385 8401 32419
rect 8435 32385 8447 32419
rect 8588 32418 8659 32446
rect 8647 32415 8659 32418
rect 8693 32415 8705 32449
rect 8647 32409 8705 32415
rect 9784 32416 9812 32524
rect 9858 32512 9864 32564
rect 9916 32552 9922 32564
rect 12986 32552 12992 32564
rect 9916 32524 12992 32552
rect 9916 32512 9922 32524
rect 12986 32512 12992 32524
rect 13044 32512 13050 32564
rect 13538 32512 13544 32564
rect 13596 32512 13602 32564
rect 11974 32444 11980 32496
rect 12032 32484 12038 32496
rect 13556 32484 13584 32512
rect 12032 32456 13584 32484
rect 12032 32444 12038 32456
rect 10318 32425 10324 32428
rect 10287 32419 10324 32425
rect 10287 32416 10299 32419
rect 9784 32388 10299 32416
rect 8389 32379 8447 32385
rect 10287 32385 10299 32388
rect 10287 32379 10324 32385
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 1854 32212 1860 32224
rect 1627 32184 1860 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 1854 32172 1860 32184
rect 1912 32172 1918 32224
rect 8018 32172 8024 32224
rect 8076 32172 8082 32224
rect 8404 32212 8432 32379
rect 10318 32376 10324 32379
rect 10376 32376 10382 32428
rect 11054 32376 11060 32428
rect 11112 32416 11118 32428
rect 11759 32419 11817 32425
rect 11759 32416 11771 32419
rect 11112 32388 11771 32416
rect 11112 32376 11118 32388
rect 11759 32385 11771 32388
rect 11805 32385 11817 32419
rect 11759 32379 11817 32385
rect 12986 32376 12992 32428
rect 13044 32376 13050 32428
rect 13541 32419 13599 32425
rect 13541 32385 13553 32419
rect 13587 32385 13599 32419
rect 13541 32379 13599 32385
rect 13909 32419 13967 32425
rect 13909 32385 13921 32419
rect 13955 32385 13967 32419
rect 13909 32379 13967 32385
rect 10045 32351 10103 32357
rect 10045 32348 10057 32351
rect 9324 32320 10057 32348
rect 9324 32212 9352 32320
rect 10045 32317 10057 32320
rect 10091 32317 10103 32351
rect 11514 32348 11520 32360
rect 10045 32311 10103 32317
rect 10980 32320 11520 32348
rect 8404 32184 9352 32212
rect 9398 32172 9404 32224
rect 9456 32172 9462 32224
rect 10060 32212 10088 32311
rect 10980 32212 11008 32320
rect 11514 32308 11520 32320
rect 11572 32308 11578 32360
rect 11057 32283 11115 32289
rect 11057 32249 11069 32283
rect 11103 32249 11115 32283
rect 13556 32280 13584 32379
rect 13924 32348 13952 32379
rect 14090 32376 14096 32428
rect 14148 32376 14154 32428
rect 14182 32348 14188 32360
rect 13924 32320 14188 32348
rect 14182 32308 14188 32320
rect 14240 32308 14246 32360
rect 11057 32243 11115 32249
rect 12406 32252 12664 32280
rect 13556 32252 14044 32280
rect 10060 32184 11008 32212
rect 11072 32212 11100 32243
rect 12406 32212 12434 32252
rect 12636 32224 12664 32252
rect 14016 32224 14044 32252
rect 11072 32184 12434 32212
rect 12526 32172 12532 32224
rect 12584 32172 12590 32224
rect 12618 32172 12624 32224
rect 12676 32172 12682 32224
rect 13265 32215 13323 32221
rect 13265 32181 13277 32215
rect 13311 32212 13323 32215
rect 13538 32212 13544 32224
rect 13311 32184 13544 32212
rect 13311 32181 13323 32184
rect 13265 32175 13323 32181
rect 13538 32172 13544 32184
rect 13596 32172 13602 32224
rect 13998 32172 14004 32224
rect 14056 32172 14062 32224
rect 14369 32215 14427 32221
rect 14369 32181 14381 32215
rect 14415 32212 14427 32215
rect 15102 32212 15108 32224
rect 14415 32184 15108 32212
rect 14415 32181 14427 32184
rect 14369 32175 14427 32181
rect 15102 32172 15108 32184
rect 15160 32172 15166 32224
rect 1104 32122 14812 32144
rect 1104 32070 2663 32122
rect 2715 32070 2727 32122
rect 2779 32070 2791 32122
rect 2843 32070 2855 32122
rect 2907 32070 2919 32122
rect 2971 32070 6090 32122
rect 6142 32070 6154 32122
rect 6206 32070 6218 32122
rect 6270 32070 6282 32122
rect 6334 32070 6346 32122
rect 6398 32070 9517 32122
rect 9569 32070 9581 32122
rect 9633 32070 9645 32122
rect 9697 32070 9709 32122
rect 9761 32070 9773 32122
rect 9825 32070 12944 32122
rect 12996 32070 13008 32122
rect 13060 32070 13072 32122
rect 13124 32070 13136 32122
rect 13188 32070 13200 32122
rect 13252 32070 14812 32122
rect 1104 32048 14812 32070
rect 6454 31968 6460 32020
rect 6512 32008 6518 32020
rect 8294 32008 8300 32020
rect 6512 31980 8300 32008
rect 6512 31968 6518 31980
rect 8294 31968 8300 31980
rect 8352 31968 8358 32020
rect 8938 31968 8944 32020
rect 8996 31968 9002 32020
rect 10410 31968 10416 32020
rect 10468 32008 10474 32020
rect 10505 32011 10563 32017
rect 10505 32008 10517 32011
rect 10468 31980 10517 32008
rect 10468 31968 10474 31980
rect 10505 31977 10517 31980
rect 10551 31977 10563 32011
rect 10505 31971 10563 31977
rect 10778 31968 10784 32020
rect 10836 31968 10842 32020
rect 11057 32011 11115 32017
rect 11057 31977 11069 32011
rect 11103 32008 11115 32011
rect 12342 32008 12348 32020
rect 11103 31980 12348 32008
rect 11103 31977 11115 31980
rect 11057 31971 11115 31977
rect 12342 31968 12348 31980
rect 12400 31968 12406 32020
rect 14093 32011 14151 32017
rect 14093 31977 14105 32011
rect 14139 32008 14151 32011
rect 14274 32008 14280 32020
rect 14139 31980 14280 32008
rect 14139 31977 14151 31980
rect 14093 31971 14151 31977
rect 14274 31968 14280 31980
rect 14332 31968 14338 32020
rect 11974 31940 11980 31952
rect 10704 31912 11980 31940
rect 6638 31872 6644 31884
rect 2746 31844 6644 31872
rect 1854 31764 1860 31816
rect 1912 31804 1918 31816
rect 2746 31804 2774 31844
rect 6638 31832 6644 31844
rect 6696 31872 6702 31884
rect 7190 31872 7196 31884
rect 6696 31844 7196 31872
rect 6696 31832 6702 31844
rect 7190 31832 7196 31844
rect 7248 31832 7254 31884
rect 1912 31776 2774 31804
rect 1912 31764 1918 31776
rect 7466 31764 7472 31816
rect 7524 31804 7530 31816
rect 10704 31813 10732 31912
rect 11974 31900 11980 31912
rect 12032 31900 12038 31952
rect 12526 31900 12532 31952
rect 12584 31940 12590 31952
rect 12584 31912 12664 31940
rect 12584 31900 12590 31912
rect 12636 31881 12664 31912
rect 13998 31900 14004 31952
rect 14056 31940 14062 31952
rect 14458 31940 14464 31952
rect 14056 31912 14464 31940
rect 14056 31900 14062 31912
rect 14458 31900 14464 31912
rect 14516 31900 14522 31952
rect 12627 31875 12685 31881
rect 12627 31841 12639 31875
rect 12673 31841 12685 31875
rect 12627 31835 12685 31841
rect 13814 31832 13820 31884
rect 13872 31832 13878 31884
rect 9125 31807 9183 31813
rect 9125 31804 9137 31807
rect 7524 31776 9137 31804
rect 7524 31764 7530 31776
rect 9125 31773 9137 31776
rect 9171 31773 9183 31807
rect 9125 31767 9183 31773
rect 10689 31807 10747 31813
rect 10689 31773 10701 31807
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 10778 31764 10784 31816
rect 10836 31804 10842 31816
rect 10965 31807 11023 31813
rect 10965 31804 10977 31807
rect 10836 31776 10977 31804
rect 10836 31764 10842 31776
rect 10965 31773 10977 31776
rect 11011 31773 11023 31807
rect 11241 31807 11299 31813
rect 11241 31804 11253 31807
rect 10965 31767 11023 31773
rect 11072 31776 11253 31804
rect 6914 31696 6920 31748
rect 6972 31736 6978 31748
rect 7190 31736 7196 31748
rect 6972 31708 7196 31736
rect 6972 31696 6978 31708
rect 7190 31696 7196 31708
rect 7248 31696 7254 31748
rect 10870 31696 10876 31748
rect 10928 31736 10934 31748
rect 11072 31736 11100 31776
rect 11241 31773 11253 31776
rect 11287 31773 11299 31807
rect 11241 31767 11299 31773
rect 11514 31764 11520 31816
rect 11572 31764 11578 31816
rect 11606 31764 11612 31816
rect 11664 31804 11670 31816
rect 11885 31807 11943 31813
rect 11885 31804 11897 31807
rect 11664 31776 11897 31804
rect 11664 31764 11670 31776
rect 11885 31773 11897 31776
rect 11931 31773 11943 31807
rect 11885 31767 11943 31773
rect 11974 31764 11980 31816
rect 12032 31764 12038 31816
rect 12161 31807 12219 31813
rect 12161 31773 12173 31807
rect 12207 31804 12219 31807
rect 12342 31804 12348 31816
rect 12207 31776 12348 31804
rect 12207 31773 12219 31776
rect 12161 31767 12219 31773
rect 12342 31764 12348 31776
rect 12400 31764 12406 31816
rect 12894 31764 12900 31816
rect 12952 31764 12958 31816
rect 13078 31813 13084 31816
rect 13035 31807 13084 31813
rect 13035 31773 13047 31807
rect 13081 31773 13084 31807
rect 13035 31767 13084 31773
rect 13078 31764 13084 31767
rect 13136 31764 13142 31816
rect 13170 31764 13176 31816
rect 13228 31764 13234 31816
rect 14274 31764 14280 31816
rect 14332 31764 14338 31816
rect 10928 31708 11100 31736
rect 11532 31708 12204 31736
rect 10928 31696 10934 31708
rect 6546 31628 6552 31680
rect 6604 31668 6610 31680
rect 9122 31668 9128 31680
rect 6604 31640 9128 31668
rect 6604 31628 6610 31640
rect 9122 31628 9128 31640
rect 9180 31628 9186 31680
rect 9306 31628 9312 31680
rect 9364 31668 9370 31680
rect 11532 31668 11560 31708
rect 9364 31640 11560 31668
rect 12176 31668 12204 31708
rect 13446 31668 13452 31680
rect 12176 31640 13452 31668
rect 9364 31628 9370 31640
rect 13446 31628 13452 31640
rect 13504 31628 13510 31680
rect 1104 31578 14971 31600
rect 1104 31526 4376 31578
rect 4428 31526 4440 31578
rect 4492 31526 4504 31578
rect 4556 31526 4568 31578
rect 4620 31526 4632 31578
rect 4684 31526 7803 31578
rect 7855 31526 7867 31578
rect 7919 31526 7931 31578
rect 7983 31526 7995 31578
rect 8047 31526 8059 31578
rect 8111 31526 11230 31578
rect 11282 31526 11294 31578
rect 11346 31526 11358 31578
rect 11410 31526 11422 31578
rect 11474 31526 11486 31578
rect 11538 31526 14657 31578
rect 14709 31526 14721 31578
rect 14773 31526 14785 31578
rect 14837 31526 14849 31578
rect 14901 31526 14913 31578
rect 14965 31526 14971 31578
rect 1104 31504 14971 31526
rect 10689 31467 10747 31473
rect 10689 31433 10701 31467
rect 10735 31464 10747 31467
rect 10778 31464 10784 31476
rect 10735 31436 10784 31464
rect 10735 31433 10747 31436
rect 10689 31427 10747 31433
rect 10778 31424 10784 31436
rect 10836 31424 10842 31476
rect 10870 31424 10876 31476
rect 10928 31464 10934 31476
rect 10965 31467 11023 31473
rect 10965 31464 10977 31467
rect 10928 31436 10977 31464
rect 10928 31424 10934 31436
rect 10965 31433 10977 31436
rect 11011 31433 11023 31467
rect 10965 31427 11023 31433
rect 11882 31424 11888 31476
rect 11940 31464 11946 31476
rect 11940 31436 13216 31464
rect 11940 31424 11946 31436
rect 6638 31356 6644 31408
rect 6696 31396 6702 31408
rect 7558 31396 7564 31408
rect 6696 31368 7564 31396
rect 6696 31356 6702 31368
rect 7558 31356 7564 31368
rect 7616 31356 7622 31408
rect 9030 31356 9036 31408
rect 9088 31396 9094 31408
rect 13188 31396 13216 31436
rect 13357 31399 13415 31405
rect 13357 31396 13369 31399
rect 9088 31368 11192 31396
rect 13188 31368 13369 31396
rect 9088 31356 9094 31368
rect 750 31288 756 31340
rect 808 31328 814 31340
rect 1397 31331 1455 31337
rect 1397 31328 1409 31331
rect 808 31300 1409 31328
rect 808 31288 814 31300
rect 1397 31297 1409 31300
rect 1443 31297 1455 31331
rect 1397 31291 1455 31297
rect 2222 31288 2228 31340
rect 2280 31328 2286 31340
rect 6822 31328 6828 31340
rect 2280 31300 6828 31328
rect 2280 31288 2286 31300
rect 6822 31288 6828 31300
rect 6880 31328 6886 31340
rect 8478 31328 8484 31340
rect 6880 31300 8484 31328
rect 6880 31288 6886 31300
rect 8478 31288 8484 31300
rect 8536 31328 8542 31340
rect 9309 31331 9367 31337
rect 9309 31328 9321 31331
rect 8536 31300 9321 31328
rect 8536 31288 8542 31300
rect 9309 31297 9321 31300
rect 9355 31297 9367 31331
rect 9309 31291 9367 31297
rect 9583 31331 9641 31337
rect 9583 31297 9595 31331
rect 9629 31328 9641 31331
rect 10134 31328 10140 31340
rect 9629 31300 10140 31328
rect 9629 31297 9641 31300
rect 9583 31291 9641 31297
rect 10134 31288 10140 31300
rect 10192 31288 10198 31340
rect 10870 31288 10876 31340
rect 10928 31288 10934 31340
rect 11164 31337 11192 31368
rect 13357 31365 13369 31368
rect 13403 31365 13415 31399
rect 13357 31359 13415 31365
rect 13446 31356 13452 31408
rect 13504 31396 13510 31408
rect 13541 31399 13599 31405
rect 13541 31396 13553 31399
rect 13504 31368 13553 31396
rect 13504 31356 13510 31368
rect 13541 31365 13553 31368
rect 13587 31365 13599 31399
rect 13541 31359 13599 31365
rect 11149 31331 11207 31337
rect 11149 31297 11161 31331
rect 11195 31297 11207 31331
rect 11701 31331 11759 31337
rect 11701 31328 11713 31331
rect 11149 31291 11207 31297
rect 11256 31300 11713 31328
rect 11256 31272 11284 31300
rect 11701 31297 11713 31300
rect 11747 31328 11759 31331
rect 11882 31328 11888 31340
rect 11747 31300 11888 31328
rect 11747 31297 11759 31300
rect 11701 31291 11759 31297
rect 11882 31288 11888 31300
rect 11940 31288 11946 31340
rect 12710 31288 12716 31340
rect 12768 31288 12774 31340
rect 14090 31288 14096 31340
rect 14148 31288 14154 31340
rect 11238 31220 11244 31272
rect 11296 31220 11302 31272
rect 11517 31263 11575 31269
rect 11517 31229 11529 31263
rect 11563 31229 11575 31263
rect 11517 31223 11575 31229
rect 11532 31192 11560 31223
rect 12158 31220 12164 31272
rect 12216 31220 12222 31272
rect 12434 31220 12440 31272
rect 12492 31220 12498 31272
rect 12526 31220 12532 31272
rect 12584 31269 12590 31272
rect 12584 31263 12612 31269
rect 12600 31229 12612 31263
rect 12584 31223 12612 31229
rect 12584 31220 12590 31223
rect 13262 31220 13268 31272
rect 13320 31260 13326 31272
rect 13630 31260 13636 31272
rect 13320 31232 13636 31260
rect 13320 31220 13326 31232
rect 13630 31220 13636 31232
rect 13688 31220 13694 31272
rect 11882 31192 11888 31204
rect 11532 31164 11888 31192
rect 11882 31152 11888 31164
rect 11940 31152 11946 31204
rect 1210 31084 1216 31136
rect 1268 31124 1274 31136
rect 1581 31127 1639 31133
rect 1581 31124 1593 31127
rect 1268 31096 1593 31124
rect 1268 31084 1274 31096
rect 1581 31093 1593 31096
rect 1627 31093 1639 31127
rect 1581 31087 1639 31093
rect 10321 31127 10379 31133
rect 10321 31093 10333 31127
rect 10367 31124 10379 31127
rect 10410 31124 10416 31136
rect 10367 31096 10416 31124
rect 10367 31093 10379 31096
rect 10321 31087 10379 31093
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10778 31084 10784 31136
rect 10836 31124 10842 31136
rect 12526 31124 12532 31136
rect 10836 31096 12532 31124
rect 10836 31084 10842 31096
rect 12526 31084 12532 31096
rect 12584 31084 12590 31136
rect 13814 31084 13820 31136
rect 13872 31084 13878 31136
rect 14369 31127 14427 31133
rect 14369 31093 14381 31127
rect 14415 31124 14427 31127
rect 15746 31124 15752 31136
rect 14415 31096 15752 31124
rect 14415 31093 14427 31096
rect 14369 31087 14427 31093
rect 15746 31084 15752 31096
rect 15804 31084 15810 31136
rect 1104 31034 14812 31056
rect 1104 30982 2663 31034
rect 2715 30982 2727 31034
rect 2779 30982 2791 31034
rect 2843 30982 2855 31034
rect 2907 30982 2919 31034
rect 2971 30982 6090 31034
rect 6142 30982 6154 31034
rect 6206 30982 6218 31034
rect 6270 30982 6282 31034
rect 6334 30982 6346 31034
rect 6398 30982 9517 31034
rect 9569 30982 9581 31034
rect 9633 30982 9645 31034
rect 9697 30982 9709 31034
rect 9761 30982 9773 31034
rect 9825 30982 12944 31034
rect 12996 30982 13008 31034
rect 13060 30982 13072 31034
rect 13124 30982 13136 31034
rect 13188 30982 13200 31034
rect 13252 30982 14812 31034
rect 1104 30960 14812 30982
rect 6730 30880 6736 30932
rect 6788 30920 6794 30932
rect 10870 30920 10876 30932
rect 6788 30892 10876 30920
rect 6788 30880 6794 30892
rect 10870 30880 10876 30892
rect 10928 30880 10934 30932
rect 13906 30880 13912 30932
rect 13964 30880 13970 30932
rect 10318 30812 10324 30864
rect 10376 30852 10382 30864
rect 10376 30824 12296 30852
rect 10376 30812 10382 30824
rect 7006 30744 7012 30796
rect 7064 30784 7070 30796
rect 7193 30787 7251 30793
rect 7193 30784 7205 30787
rect 7064 30756 7205 30784
rect 7064 30744 7070 30756
rect 7193 30753 7205 30756
rect 7239 30753 7251 30787
rect 7193 30747 7251 30753
rect 1394 30676 1400 30728
rect 1452 30676 1458 30728
rect 7208 30716 7236 30747
rect 8662 30744 8668 30796
rect 8720 30784 8726 30796
rect 8846 30784 8852 30796
rect 8720 30756 8852 30784
rect 8720 30744 8726 30756
rect 8846 30744 8852 30756
rect 8904 30744 8910 30796
rect 11333 30787 11391 30793
rect 11333 30753 11345 30787
rect 11379 30784 11391 30787
rect 11790 30784 11796 30796
rect 11379 30756 11796 30784
rect 11379 30753 11391 30756
rect 11333 30747 11391 30753
rect 11790 30744 11796 30756
rect 11848 30744 11854 30796
rect 7208 30688 7328 30716
rect 7300 30592 7328 30688
rect 7451 30689 7509 30695
rect 7451 30655 7463 30689
rect 7497 30686 7509 30689
rect 7497 30655 7512 30686
rect 10502 30676 10508 30728
rect 10560 30716 10566 30728
rect 12268 30725 12296 30824
rect 12710 30812 12716 30864
rect 12768 30812 12774 30864
rect 12618 30744 12624 30796
rect 12676 30784 12682 30796
rect 12802 30784 12808 30796
rect 12676 30756 12808 30784
rect 12676 30744 12682 30756
rect 12802 30744 12808 30756
rect 12860 30784 12866 30796
rect 12989 30787 13047 30793
rect 12989 30784 13001 30787
rect 12860 30756 13001 30784
rect 12860 30744 12866 30756
rect 12989 30753 13001 30756
rect 13035 30753 13047 30787
rect 12989 30747 13047 30753
rect 13265 30787 13323 30793
rect 13265 30753 13277 30787
rect 13311 30784 13323 30787
rect 13630 30784 13636 30796
rect 13311 30756 13636 30784
rect 13311 30753 13323 30756
rect 13265 30747 13323 30753
rect 13630 30744 13636 30756
rect 13688 30744 13694 30796
rect 13170 30725 13176 30728
rect 11609 30719 11667 30725
rect 11609 30716 11621 30719
rect 10560 30688 11621 30716
rect 10560 30676 10566 30688
rect 11609 30685 11621 30688
rect 11655 30685 11667 30719
rect 11609 30679 11667 30685
rect 12069 30719 12127 30725
rect 12069 30685 12081 30719
rect 12115 30685 12127 30719
rect 12069 30679 12127 30685
rect 12253 30719 12311 30725
rect 12253 30685 12265 30719
rect 12299 30685 12311 30719
rect 12253 30679 12311 30685
rect 13127 30719 13176 30725
rect 13127 30685 13139 30719
rect 13173 30685 13176 30719
rect 13127 30679 13176 30685
rect 7451 30649 7512 30655
rect 7484 30648 7512 30649
rect 7484 30620 8708 30648
rect 8680 30592 8708 30620
rect 11054 30608 11060 30660
rect 11112 30608 11118 30660
rect 11974 30608 11980 30660
rect 12032 30608 12038 30660
rect 12084 30648 12112 30679
rect 13170 30676 13176 30679
rect 13228 30676 13234 30728
rect 12084 30620 12296 30648
rect 1581 30583 1639 30589
rect 1581 30549 1593 30583
rect 1627 30580 1639 30583
rect 5258 30580 5264 30592
rect 1627 30552 5264 30580
rect 1627 30549 1639 30552
rect 1581 30543 1639 30549
rect 5258 30540 5264 30552
rect 5316 30540 5322 30592
rect 7282 30540 7288 30592
rect 7340 30540 7346 30592
rect 8205 30583 8263 30589
rect 8205 30549 8217 30583
rect 8251 30580 8263 30583
rect 8386 30580 8392 30592
rect 8251 30552 8392 30580
rect 8251 30549 8263 30552
rect 8205 30543 8263 30549
rect 8386 30540 8392 30552
rect 8444 30540 8450 30592
rect 8662 30540 8668 30592
rect 8720 30540 8726 30592
rect 10134 30540 10140 30592
rect 10192 30580 10198 30592
rect 12066 30580 12072 30592
rect 10192 30552 12072 30580
rect 10192 30540 10198 30552
rect 12066 30540 12072 30552
rect 12124 30540 12130 30592
rect 12268 30580 12296 30620
rect 12434 30580 12440 30592
rect 12268 30552 12440 30580
rect 12434 30540 12440 30552
rect 12492 30540 12498 30592
rect 1104 30490 14971 30512
rect 1104 30438 4376 30490
rect 4428 30438 4440 30490
rect 4492 30438 4504 30490
rect 4556 30438 4568 30490
rect 4620 30438 4632 30490
rect 4684 30438 7803 30490
rect 7855 30438 7867 30490
rect 7919 30438 7931 30490
rect 7983 30438 7995 30490
rect 8047 30438 8059 30490
rect 8111 30438 11230 30490
rect 11282 30438 11294 30490
rect 11346 30438 11358 30490
rect 11410 30438 11422 30490
rect 11474 30438 11486 30490
rect 11538 30438 14657 30490
rect 14709 30438 14721 30490
rect 14773 30438 14785 30490
rect 14837 30438 14849 30490
rect 14901 30438 14913 30490
rect 14965 30438 14971 30490
rect 1104 30416 14971 30438
rect 6638 30336 6644 30388
rect 6696 30376 6702 30388
rect 8570 30376 8576 30388
rect 6696 30348 8576 30376
rect 6696 30336 6702 30348
rect 8570 30336 8576 30348
rect 8628 30336 8634 30388
rect 9306 30336 9312 30388
rect 9364 30376 9370 30388
rect 9490 30376 9496 30388
rect 9364 30348 9496 30376
rect 9364 30336 9370 30348
rect 9490 30336 9496 30348
rect 9548 30336 9554 30388
rect 10870 30336 10876 30388
rect 10928 30376 10934 30388
rect 10928 30348 11100 30376
rect 10928 30336 10934 30348
rect 7466 30268 7472 30320
rect 7524 30268 7530 30320
rect 10045 30311 10103 30317
rect 10045 30277 10057 30311
rect 10091 30308 10103 30311
rect 10965 30311 11023 30317
rect 10965 30308 10977 30311
rect 10091 30280 10977 30308
rect 10091 30277 10103 30280
rect 10045 30271 10103 30277
rect 10965 30277 10977 30280
rect 11011 30277 11023 30311
rect 10965 30271 11023 30277
rect 6546 30200 6552 30252
rect 6604 30240 6610 30252
rect 6825 30243 6883 30249
rect 6825 30240 6837 30243
rect 6604 30212 6837 30240
rect 6604 30200 6610 30212
rect 6825 30209 6837 30212
rect 6871 30209 6883 30243
rect 6825 30203 6883 30209
rect 6840 30036 6868 30203
rect 7006 30200 7012 30252
rect 7064 30240 7070 30252
rect 7099 30243 7157 30249
rect 7099 30240 7111 30243
rect 7064 30212 7111 30240
rect 7064 30200 7070 30212
rect 7099 30209 7111 30212
rect 7145 30240 7157 30243
rect 7484 30240 7512 30268
rect 7145 30212 7512 30240
rect 7145 30209 7157 30212
rect 7099 30203 7157 30209
rect 9398 30200 9404 30252
rect 9456 30200 9462 30252
rect 10413 30243 10471 30249
rect 10413 30209 10425 30243
rect 10459 30240 10471 30243
rect 10870 30240 10876 30252
rect 10459 30212 10876 30240
rect 10459 30209 10471 30212
rect 10413 30203 10471 30209
rect 10870 30200 10876 30212
rect 10928 30200 10934 30252
rect 11072 30240 11100 30348
rect 11330 30268 11336 30320
rect 11388 30268 11394 30320
rect 11514 30240 11520 30252
rect 11072 30212 11520 30240
rect 11514 30200 11520 30212
rect 11572 30200 11578 30252
rect 11793 30243 11851 30249
rect 11793 30209 11805 30243
rect 11839 30209 11851 30243
rect 11793 30203 11851 30209
rect 12159 30243 12217 30249
rect 12159 30209 12171 30243
rect 12205 30240 12217 30243
rect 12250 30240 12256 30252
rect 12205 30212 12256 30240
rect 12205 30209 12217 30212
rect 12159 30203 12217 30209
rect 8110 30132 8116 30184
rect 8168 30172 8174 30184
rect 8205 30175 8263 30181
rect 8205 30172 8217 30175
rect 8168 30144 8217 30172
rect 8168 30132 8174 30144
rect 8205 30141 8217 30144
rect 8251 30141 8263 30175
rect 8205 30135 8263 30141
rect 8389 30175 8447 30181
rect 8389 30141 8401 30175
rect 8435 30172 8447 30175
rect 8478 30172 8484 30184
rect 8435 30144 8484 30172
rect 8435 30141 8447 30144
rect 8389 30135 8447 30141
rect 8478 30132 8484 30144
rect 8536 30132 8542 30184
rect 9306 30181 9312 30184
rect 9125 30175 9183 30181
rect 9125 30172 9137 30175
rect 8956 30144 9137 30172
rect 8956 30116 8984 30144
rect 9125 30141 9137 30144
rect 9171 30141 9183 30175
rect 9125 30135 9183 30141
rect 9263 30175 9312 30181
rect 9263 30141 9275 30175
rect 9309 30141 9312 30175
rect 9263 30135 9312 30141
rect 9306 30132 9312 30135
rect 9364 30132 9370 30184
rect 10134 30132 10140 30184
rect 10192 30172 10198 30184
rect 11808 30172 11836 30203
rect 12250 30200 12256 30212
rect 12308 30200 12314 30252
rect 13541 30243 13599 30249
rect 13541 30209 13553 30243
rect 13587 30209 13599 30243
rect 13541 30203 13599 30209
rect 13909 30243 13967 30249
rect 13909 30209 13921 30243
rect 13955 30209 13967 30243
rect 13909 30203 13967 30209
rect 14093 30243 14151 30249
rect 14093 30209 14105 30243
rect 14139 30240 14151 30243
rect 15562 30240 15568 30252
rect 14139 30212 15568 30240
rect 14139 30209 14151 30212
rect 14093 30203 14151 30209
rect 10192 30144 11836 30172
rect 11885 30175 11943 30181
rect 10192 30132 10198 30144
rect 11885 30141 11897 30175
rect 11931 30141 11943 30175
rect 11885 30135 11943 30141
rect 7837 30107 7895 30113
rect 7837 30073 7849 30107
rect 7883 30104 7895 30107
rect 8849 30107 8907 30113
rect 8849 30104 8861 30107
rect 7883 30076 8861 30104
rect 7883 30073 7895 30076
rect 7837 30067 7895 30073
rect 8849 30073 8861 30076
rect 8895 30073 8907 30107
rect 8849 30067 8907 30073
rect 8938 30064 8944 30116
rect 8996 30064 9002 30116
rect 11146 30064 11152 30116
rect 11204 30104 11210 30116
rect 11609 30107 11667 30113
rect 11609 30104 11621 30107
rect 11204 30076 11621 30104
rect 11204 30064 11210 30076
rect 11609 30073 11621 30076
rect 11655 30073 11667 30107
rect 11609 30067 11667 30073
rect 7282 30036 7288 30048
rect 6840 30008 7288 30036
rect 7282 29996 7288 30008
rect 7340 30036 7346 30048
rect 9950 30036 9956 30048
rect 7340 30008 9956 30036
rect 7340 29996 7346 30008
rect 9950 29996 9956 30008
rect 10008 29996 10014 30048
rect 10689 30039 10747 30045
rect 10689 30005 10701 30039
rect 10735 30036 10747 30039
rect 10962 30036 10968 30048
rect 10735 30008 10968 30036
rect 10735 30005 10747 30008
rect 10689 29999 10747 30005
rect 10962 29996 10968 30008
rect 11020 29996 11026 30048
rect 11238 29996 11244 30048
rect 11296 30036 11302 30048
rect 11900 30036 11928 30135
rect 13556 30104 13584 30203
rect 13924 30172 13952 30203
rect 15562 30200 15568 30212
rect 15620 30200 15626 30252
rect 15470 30172 15476 30184
rect 13924 30144 15476 30172
rect 15470 30132 15476 30144
rect 15528 30132 15534 30184
rect 13906 30104 13912 30116
rect 13556 30076 13912 30104
rect 13906 30064 13912 30076
rect 13964 30064 13970 30116
rect 11296 30008 11928 30036
rect 11296 29996 11302 30008
rect 12158 29996 12164 30048
rect 12216 30036 12222 30048
rect 12618 30036 12624 30048
rect 12216 30008 12624 30036
rect 12216 29996 12222 30008
rect 12618 29996 12624 30008
rect 12676 29996 12682 30048
rect 12894 29996 12900 30048
rect 12952 29996 12958 30048
rect 14369 30039 14427 30045
rect 14369 30005 14381 30039
rect 14415 30036 14427 30039
rect 14550 30036 14556 30048
rect 14415 30008 14556 30036
rect 14415 30005 14427 30008
rect 14369 29999 14427 30005
rect 14550 29996 14556 30008
rect 14608 29996 14614 30048
rect 15102 29996 15108 30048
rect 15160 30036 15166 30048
rect 15562 30036 15568 30048
rect 15160 30008 15568 30036
rect 15160 29996 15166 30008
rect 15562 29996 15568 30008
rect 15620 29996 15626 30048
rect 1104 29946 14812 29968
rect 1104 29894 2663 29946
rect 2715 29894 2727 29946
rect 2779 29894 2791 29946
rect 2843 29894 2855 29946
rect 2907 29894 2919 29946
rect 2971 29894 6090 29946
rect 6142 29894 6154 29946
rect 6206 29894 6218 29946
rect 6270 29894 6282 29946
rect 6334 29894 6346 29946
rect 6398 29894 9517 29946
rect 9569 29894 9581 29946
rect 9633 29894 9645 29946
rect 9697 29894 9709 29946
rect 9761 29894 9773 29946
rect 9825 29894 12944 29946
rect 12996 29894 13008 29946
rect 13060 29894 13072 29946
rect 13124 29894 13136 29946
rect 13188 29894 13200 29946
rect 13252 29894 14812 29946
rect 1104 29872 14812 29894
rect 8110 29792 8116 29844
rect 8168 29832 8174 29844
rect 10042 29832 10048 29844
rect 8168 29804 10048 29832
rect 8168 29792 8174 29804
rect 10042 29792 10048 29804
rect 10100 29792 10106 29844
rect 10686 29832 10692 29844
rect 10336 29804 10692 29832
rect 9950 29724 9956 29776
rect 10008 29764 10014 29776
rect 10336 29764 10364 29804
rect 10686 29792 10692 29804
rect 10744 29792 10750 29844
rect 10778 29792 10784 29844
rect 10836 29832 10842 29844
rect 10836 29804 12388 29832
rect 10836 29792 10842 29804
rect 10008 29736 10364 29764
rect 10008 29724 10014 29736
rect 8570 29656 8576 29708
rect 8628 29696 8634 29708
rect 8941 29699 8999 29705
rect 8941 29696 8953 29699
rect 8628 29668 8953 29696
rect 8628 29656 8634 29668
rect 8941 29665 8953 29668
rect 8987 29665 8999 29699
rect 8941 29659 8999 29665
rect 750 29588 756 29640
rect 808 29628 814 29640
rect 1397 29631 1455 29637
rect 1397 29628 1409 29631
rect 808 29600 1409 29628
rect 808 29588 814 29600
rect 1397 29597 1409 29600
rect 1443 29597 1455 29631
rect 10134 29628 10140 29640
rect 1397 29591 1455 29597
rect 9215 29621 9273 29627
rect 9215 29587 9227 29621
rect 9261 29618 9273 29621
rect 9324 29618 10140 29628
rect 9261 29600 10140 29618
rect 9261 29590 9352 29600
rect 9261 29587 9273 29590
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 10336 29637 10364 29736
rect 11330 29724 11336 29776
rect 11388 29724 11394 29776
rect 12360 29764 12388 29804
rect 12618 29792 12624 29844
rect 12676 29832 12682 29844
rect 12713 29835 12771 29841
rect 12713 29832 12725 29835
rect 12676 29804 12725 29832
rect 12676 29792 12682 29804
rect 12713 29801 12725 29804
rect 12759 29801 12771 29835
rect 12713 29795 12771 29801
rect 13538 29764 13544 29776
rect 12360 29736 13544 29764
rect 13538 29724 13544 29736
rect 13596 29724 13602 29776
rect 12618 29696 12624 29708
rect 12314 29668 12624 29696
rect 10321 29631 10379 29637
rect 10321 29597 10333 29631
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 10595 29631 10653 29637
rect 10595 29597 10607 29631
rect 10641 29628 10653 29631
rect 11238 29628 11244 29640
rect 10641 29600 11244 29628
rect 10641 29597 10653 29600
rect 10595 29591 10653 29597
rect 11238 29588 11244 29600
rect 11296 29588 11302 29640
rect 11422 29588 11428 29640
rect 11480 29628 11486 29640
rect 11701 29631 11759 29637
rect 11701 29628 11713 29631
rect 11480 29600 11713 29628
rect 11480 29588 11486 29600
rect 11701 29597 11713 29600
rect 11747 29597 11759 29631
rect 11701 29591 11759 29597
rect 11975 29631 12033 29637
rect 11975 29597 11987 29631
rect 12021 29628 12033 29631
rect 12314 29628 12342 29668
rect 12618 29656 12624 29668
rect 12676 29696 12682 29708
rect 12676 29668 13768 29696
rect 12676 29656 12682 29668
rect 13740 29640 13768 29668
rect 12021 29600 12342 29628
rect 12021 29597 12033 29600
rect 11975 29591 12033 29597
rect 13722 29588 13728 29640
rect 13780 29588 13786 29640
rect 9215 29581 9273 29587
rect 8570 29520 8576 29572
rect 8628 29560 8634 29572
rect 8628 29532 8892 29560
rect 8628 29520 8634 29532
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 1762 29492 1768 29504
rect 1627 29464 1768 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 1762 29452 1768 29464
rect 1820 29492 1826 29504
rect 8754 29492 8760 29504
rect 1820 29464 8760 29492
rect 1820 29452 1826 29464
rect 8754 29452 8760 29464
rect 8812 29452 8818 29504
rect 8864 29492 8892 29532
rect 9646 29532 10548 29560
rect 9646 29492 9674 29532
rect 8864 29464 9674 29492
rect 9950 29452 9956 29504
rect 10008 29452 10014 29504
rect 10520 29492 10548 29532
rect 11330 29520 11336 29572
rect 11388 29560 11394 29572
rect 12986 29560 12992 29572
rect 11388 29532 12992 29560
rect 11388 29520 11394 29532
rect 12986 29520 12992 29532
rect 13044 29520 13050 29572
rect 13538 29520 13544 29572
rect 13596 29520 13602 29572
rect 12618 29492 12624 29504
rect 10520 29464 12624 29492
rect 12618 29452 12624 29464
rect 12676 29452 12682 29504
rect 13630 29452 13636 29504
rect 13688 29452 13694 29504
rect 1104 29402 14971 29424
rect 1104 29350 4376 29402
rect 4428 29350 4440 29402
rect 4492 29350 4504 29402
rect 4556 29350 4568 29402
rect 4620 29350 4632 29402
rect 4684 29350 7803 29402
rect 7855 29350 7867 29402
rect 7919 29350 7931 29402
rect 7983 29350 7995 29402
rect 8047 29350 8059 29402
rect 8111 29350 11230 29402
rect 11282 29350 11294 29402
rect 11346 29350 11358 29402
rect 11410 29350 11422 29402
rect 11474 29350 11486 29402
rect 11538 29350 14657 29402
rect 14709 29350 14721 29402
rect 14773 29350 14785 29402
rect 14837 29350 14849 29402
rect 14901 29350 14913 29402
rect 14965 29350 14971 29402
rect 1104 29328 14971 29350
rect 8478 29288 8484 29300
rect 8220 29260 8484 29288
rect 1394 29112 1400 29164
rect 1452 29112 1458 29164
rect 2406 29112 2412 29164
rect 2464 29152 2470 29164
rect 8220 29161 8248 29260
rect 8478 29248 8484 29260
rect 8536 29248 8542 29300
rect 8754 29248 8760 29300
rect 8812 29288 8818 29300
rect 8812 29260 9812 29288
rect 8812 29248 8818 29260
rect 9784 29220 9812 29260
rect 9858 29248 9864 29300
rect 9916 29248 9922 29300
rect 11238 29288 11244 29300
rect 10244 29260 11244 29288
rect 10244 29220 10272 29260
rect 11238 29248 11244 29260
rect 11296 29248 11302 29300
rect 12250 29288 12256 29300
rect 11624 29260 12256 29288
rect 9784 29192 10272 29220
rect 11054 29180 11060 29232
rect 11112 29220 11118 29232
rect 11517 29223 11575 29229
rect 11517 29220 11529 29223
rect 11112 29192 11529 29220
rect 11112 29180 11118 29192
rect 11517 29189 11529 29192
rect 11563 29189 11575 29223
rect 11517 29183 11575 29189
rect 10319 29165 10377 29171
rect 8205 29155 8263 29161
rect 8205 29152 8217 29155
rect 2464 29124 8217 29152
rect 2464 29112 2470 29124
rect 8205 29121 8217 29124
rect 8251 29121 8263 29155
rect 8205 29115 8263 29121
rect 9214 29112 9220 29164
rect 9272 29112 9278 29164
rect 10319 29131 10331 29165
rect 10365 29152 10377 29165
rect 11624 29152 11652 29260
rect 12250 29248 12256 29260
rect 12308 29248 12314 29300
rect 12618 29248 12624 29300
rect 12676 29288 12682 29300
rect 12676 29260 13952 29288
rect 12676 29248 12682 29260
rect 13924 29229 13952 29260
rect 13909 29223 13967 29229
rect 13909 29189 13921 29223
rect 13955 29189 13967 29223
rect 13909 29183 13967 29189
rect 10365 29131 10916 29152
rect 10319 29125 10916 29131
rect 10336 29124 10916 29125
rect 7006 29044 7012 29096
rect 7064 29084 7070 29096
rect 8021 29087 8079 29093
rect 8021 29084 8033 29087
rect 7064 29056 8033 29084
rect 7064 29044 7070 29056
rect 8021 29053 8033 29056
rect 8067 29053 8079 29087
rect 8021 29047 8079 29053
rect 8386 29044 8392 29096
rect 8444 29084 8450 29096
rect 8665 29087 8723 29093
rect 8665 29084 8677 29087
rect 8444 29056 8677 29084
rect 8444 29044 8450 29056
rect 8665 29053 8677 29056
rect 8711 29053 8723 29087
rect 8938 29084 8944 29096
rect 8665 29047 8723 29053
rect 8772 29056 8944 29084
rect 1581 29019 1639 29025
rect 1581 28985 1593 29019
rect 1627 29016 1639 29019
rect 1946 29016 1952 29028
rect 1627 28988 1952 29016
rect 1627 28985 1639 28988
rect 1581 28979 1639 28985
rect 1946 28976 1952 28988
rect 2004 28976 2010 29028
rect 7282 28976 7288 29028
rect 7340 29016 7346 29028
rect 8772 29016 8800 29056
rect 8938 29044 8944 29056
rect 8996 29044 9002 29096
rect 9079 29087 9137 29093
rect 9079 29053 9091 29087
rect 9125 29084 9137 29087
rect 9125 29056 9628 29084
rect 9125 29053 9137 29056
rect 9079 29047 9137 29053
rect 7340 28988 8800 29016
rect 7340 28976 7346 28988
rect 8202 28908 8208 28960
rect 8260 28948 8266 28960
rect 9600 28948 9628 29056
rect 9858 29044 9864 29096
rect 9916 29084 9922 29096
rect 10045 29087 10103 29093
rect 10045 29084 10057 29087
rect 9916 29056 10057 29084
rect 9916 29044 9922 29056
rect 10045 29053 10057 29056
rect 10091 29053 10103 29087
rect 10888 29084 10916 29124
rect 11440 29124 11652 29152
rect 11440 29084 11468 29124
rect 12156 29112 12162 29164
rect 12214 29152 12220 29164
rect 13725 29155 13783 29161
rect 12214 29124 12259 29152
rect 12214 29112 12220 29124
rect 13725 29121 13737 29155
rect 13771 29152 13783 29155
rect 14182 29152 14188 29164
rect 13771 29124 14188 29152
rect 13771 29121 13783 29124
rect 13725 29115 13783 29121
rect 12299 29087 12357 29093
rect 12299 29084 12311 29087
rect 10888 29056 11468 29084
rect 11532 29056 12311 29084
rect 10045 29047 10103 29053
rect 11532 29028 11560 29056
rect 12299 29053 12311 29056
rect 12345 29053 12357 29087
rect 12299 29047 12357 29053
rect 12437 29087 12495 29093
rect 12437 29053 12449 29087
rect 12483 29084 12495 29087
rect 12713 29087 12771 29093
rect 12483 29056 12664 29084
rect 12483 29053 12495 29056
rect 12437 29047 12495 29053
rect 11238 28976 11244 29028
rect 11296 28976 11302 29028
rect 11514 28976 11520 29028
rect 11572 28976 11578 29028
rect 8260 28920 9628 28948
rect 8260 28908 8266 28920
rect 11054 28908 11060 28960
rect 11112 28908 11118 28960
rect 11256 28948 11284 28976
rect 12250 28948 12256 28960
rect 11256 28920 12256 28948
rect 12250 28908 12256 28920
rect 12308 28908 12314 28960
rect 12636 28948 12664 29056
rect 12713 29053 12725 29087
rect 12759 29084 12771 29087
rect 12986 29084 12992 29096
rect 12759 29056 12992 29084
rect 12759 29053 12771 29056
rect 12713 29047 12771 29053
rect 12986 29044 12992 29056
rect 13044 29044 13050 29096
rect 13170 29044 13176 29096
rect 13228 29044 13234 29096
rect 13357 29087 13415 29093
rect 13357 29053 13369 29087
rect 13403 29084 13415 29087
rect 13740 29084 13768 29115
rect 14182 29112 14188 29124
rect 14240 29112 14246 29164
rect 13403 29056 13768 29084
rect 13403 29053 13415 29056
rect 13357 29047 13415 29053
rect 13188 29016 13216 29044
rect 14185 29019 14243 29025
rect 13188 28988 13584 29016
rect 13556 28960 13584 28988
rect 14185 28985 14197 29019
rect 14231 29016 14243 29019
rect 15102 29016 15108 29028
rect 14231 28988 15108 29016
rect 14231 28985 14243 28988
rect 14185 28979 14243 28985
rect 15102 28976 15108 28988
rect 15160 28976 15166 29028
rect 12710 28948 12716 28960
rect 12636 28920 12716 28948
rect 12710 28908 12716 28920
rect 12768 28908 12774 28960
rect 13538 28908 13544 28960
rect 13596 28908 13602 28960
rect 1104 28858 14812 28880
rect 1104 28806 2663 28858
rect 2715 28806 2727 28858
rect 2779 28806 2791 28858
rect 2843 28806 2855 28858
rect 2907 28806 2919 28858
rect 2971 28806 6090 28858
rect 6142 28806 6154 28858
rect 6206 28806 6218 28858
rect 6270 28806 6282 28858
rect 6334 28806 6346 28858
rect 6398 28806 9517 28858
rect 9569 28806 9581 28858
rect 9633 28806 9645 28858
rect 9697 28806 9709 28858
rect 9761 28806 9773 28858
rect 9825 28806 12944 28858
rect 12996 28806 13008 28858
rect 13060 28806 13072 28858
rect 13124 28806 13136 28858
rect 13188 28806 13200 28858
rect 13252 28806 14812 28858
rect 1104 28784 14812 28806
rect 6822 28744 6828 28756
rect 6380 28716 6828 28744
rect 6380 28617 6408 28716
rect 6822 28704 6828 28716
rect 6880 28704 6886 28756
rect 7374 28704 7380 28756
rect 7432 28744 7438 28756
rect 8754 28744 8760 28756
rect 7432 28716 8760 28744
rect 7432 28704 7438 28716
rect 8754 28704 8760 28716
rect 8812 28704 8818 28756
rect 9048 28716 9444 28744
rect 6365 28611 6423 28617
rect 6365 28577 6377 28611
rect 6411 28577 6423 28611
rect 6365 28571 6423 28577
rect 9048 28552 9076 28716
rect 9306 28636 9312 28688
rect 9364 28636 9370 28688
rect 1210 28500 1216 28552
rect 1268 28540 1274 28552
rect 6638 28540 6644 28552
rect 1268 28512 2774 28540
rect 1268 28500 1274 28512
rect 2746 28472 2774 28512
rect 6472 28512 6644 28540
rect 6472 28472 6500 28512
rect 6638 28500 6644 28512
rect 6696 28500 6702 28552
rect 9030 28500 9036 28552
rect 9088 28500 9094 28552
rect 9217 28543 9275 28549
rect 9217 28509 9229 28543
rect 9263 28540 9275 28543
rect 9324 28540 9352 28636
rect 9416 28617 9444 28716
rect 9582 28704 9588 28756
rect 9640 28744 9646 28756
rect 10318 28744 10324 28756
rect 9640 28716 10324 28744
rect 9640 28704 9646 28716
rect 10318 28704 10324 28716
rect 10376 28704 10382 28756
rect 11057 28747 11115 28753
rect 11057 28713 11069 28747
rect 11103 28744 11115 28747
rect 13722 28744 13728 28756
rect 11103 28716 13728 28744
rect 11103 28713 11115 28716
rect 11057 28707 11115 28713
rect 13722 28704 13728 28716
rect 13780 28704 13786 28756
rect 13909 28747 13967 28753
rect 13909 28713 13921 28747
rect 13955 28744 13967 28747
rect 13998 28744 14004 28756
rect 13955 28716 14004 28744
rect 13955 28713 13967 28716
rect 13909 28707 13967 28713
rect 13998 28704 14004 28716
rect 14056 28704 14062 28756
rect 9861 28679 9919 28685
rect 9861 28645 9873 28679
rect 9907 28676 9919 28679
rect 9950 28676 9956 28688
rect 9907 28648 9956 28676
rect 9907 28645 9919 28648
rect 9861 28639 9919 28645
rect 9950 28636 9956 28648
rect 10008 28636 10014 28688
rect 12618 28676 12624 28688
rect 12268 28648 12624 28676
rect 9401 28611 9459 28617
rect 9401 28577 9413 28611
rect 9447 28577 9459 28611
rect 9401 28571 9459 28577
rect 9490 28568 9496 28620
rect 9548 28608 9554 28620
rect 10137 28611 10195 28617
rect 10137 28608 10149 28611
rect 9548 28580 10149 28608
rect 9548 28568 9554 28580
rect 10137 28577 10149 28580
rect 10183 28577 10195 28611
rect 10137 28571 10195 28577
rect 10410 28568 10416 28620
rect 10468 28568 10474 28620
rect 12268 28617 12296 28648
rect 12618 28636 12624 28648
rect 12676 28636 12682 28688
rect 12713 28679 12771 28685
rect 12713 28645 12725 28679
rect 12759 28676 12771 28679
rect 12802 28676 12808 28688
rect 12759 28648 12808 28676
rect 12759 28645 12771 28648
rect 12713 28639 12771 28645
rect 12802 28636 12808 28648
rect 12860 28636 12866 28688
rect 13170 28617 13176 28620
rect 12253 28611 12311 28617
rect 12253 28577 12265 28611
rect 12299 28577 12311 28611
rect 12253 28571 12311 28577
rect 13127 28611 13176 28617
rect 13127 28577 13139 28611
rect 13173 28577 13176 28611
rect 13127 28571 13176 28577
rect 13170 28568 13176 28571
rect 13228 28568 13234 28620
rect 13265 28611 13323 28617
rect 13265 28577 13277 28611
rect 13311 28608 13323 28611
rect 13814 28608 13820 28620
rect 13311 28580 13820 28608
rect 13311 28577 13323 28580
rect 13265 28571 13323 28577
rect 13814 28568 13820 28580
rect 13872 28568 13878 28620
rect 9582 28540 9588 28552
rect 9263 28512 9588 28540
rect 9263 28509 9275 28512
rect 9217 28503 9275 28509
rect 9582 28500 9588 28512
rect 9640 28500 9646 28552
rect 10318 28549 10324 28552
rect 10275 28543 10324 28549
rect 10275 28509 10287 28543
rect 10321 28509 10324 28543
rect 10275 28503 10324 28509
rect 10318 28500 10324 28503
rect 10376 28500 10382 28552
rect 12066 28500 12072 28552
rect 12124 28500 12130 28552
rect 12986 28500 12992 28552
rect 13044 28500 13050 28552
rect 2746 28444 6500 28472
rect 11609 28475 11667 28481
rect 11609 28441 11621 28475
rect 11655 28472 11667 28475
rect 11655 28444 12020 28472
rect 11655 28441 11667 28444
rect 11609 28435 11667 28441
rect 7377 28407 7435 28413
rect 7377 28373 7389 28407
rect 7423 28404 7435 28407
rect 7466 28404 7472 28416
rect 7423 28376 7472 28404
rect 7423 28373 7435 28376
rect 7377 28367 7435 28373
rect 7466 28364 7472 28376
rect 7524 28364 7530 28416
rect 10686 28364 10692 28416
rect 10744 28404 10750 28416
rect 11514 28404 11520 28416
rect 10744 28376 11520 28404
rect 10744 28364 10750 28376
rect 11514 28364 11520 28376
rect 11572 28364 11578 28416
rect 11882 28364 11888 28416
rect 11940 28364 11946 28416
rect 11992 28404 12020 28444
rect 13354 28404 13360 28416
rect 11992 28376 13360 28404
rect 13354 28364 13360 28376
rect 13412 28364 13418 28416
rect 1104 28314 14971 28336
rect 1104 28262 4376 28314
rect 4428 28262 4440 28314
rect 4492 28262 4504 28314
rect 4556 28262 4568 28314
rect 4620 28262 4632 28314
rect 4684 28262 7803 28314
rect 7855 28262 7867 28314
rect 7919 28262 7931 28314
rect 7983 28262 7995 28314
rect 8047 28262 8059 28314
rect 8111 28262 11230 28314
rect 11282 28262 11294 28314
rect 11346 28262 11358 28314
rect 11410 28262 11422 28314
rect 11474 28262 11486 28314
rect 11538 28262 14657 28314
rect 14709 28262 14721 28314
rect 14773 28262 14785 28314
rect 14837 28262 14849 28314
rect 14901 28262 14913 28314
rect 14965 28262 14971 28314
rect 1104 28240 14971 28262
rect 1394 28160 1400 28212
rect 1452 28200 1458 28212
rect 1581 28203 1639 28209
rect 1581 28200 1593 28203
rect 1452 28172 1593 28200
rect 1452 28160 1458 28172
rect 1581 28169 1593 28172
rect 1627 28200 1639 28203
rect 7374 28200 7380 28212
rect 1627 28172 7380 28200
rect 1627 28169 1639 28172
rect 1581 28163 1639 28169
rect 7374 28160 7380 28172
rect 7432 28160 7438 28212
rect 9582 28200 9588 28212
rect 8680 28172 9588 28200
rect 7558 28103 7564 28144
rect 7543 28097 7564 28103
rect 750 28024 756 28076
rect 808 28064 814 28076
rect 1397 28067 1455 28073
rect 1397 28064 1409 28067
rect 808 28036 1409 28064
rect 808 28024 814 28036
rect 1397 28033 1409 28036
rect 1443 28033 1455 28067
rect 1397 28027 1455 28033
rect 6822 28024 6828 28076
rect 6880 28064 6886 28076
rect 7285 28067 7343 28073
rect 7285 28064 7297 28067
rect 6880 28036 7297 28064
rect 6880 28024 6886 28036
rect 7285 28033 7297 28036
rect 7331 28033 7343 28067
rect 7543 28063 7555 28097
rect 7616 28092 7622 28144
rect 7589 28066 7604 28092
rect 8680 28073 8708 28172
rect 9582 28160 9588 28172
rect 9640 28160 9646 28212
rect 9950 28160 9956 28212
rect 10008 28200 10014 28212
rect 10318 28200 10324 28212
rect 10008 28172 10324 28200
rect 10008 28160 10014 28172
rect 10318 28160 10324 28172
rect 10376 28160 10382 28212
rect 10502 28160 10508 28212
rect 10560 28160 10566 28212
rect 12250 28160 12256 28212
rect 12308 28200 12314 28212
rect 12308 28172 13474 28200
rect 12308 28160 12314 28172
rect 13446 28132 13474 28172
rect 13814 28132 13820 28144
rect 13446 28104 13820 28132
rect 9766 28073 9772 28076
rect 8665 28067 8723 28073
rect 7589 28063 7601 28066
rect 7543 28057 7601 28063
rect 7285 28027 7343 28033
rect 8665 28033 8677 28067
rect 8711 28033 8723 28067
rect 8665 28027 8723 28033
rect 9723 28067 9772 28073
rect 9723 28033 9735 28067
rect 9769 28033 9772 28067
rect 9723 28027 9772 28033
rect 7098 27820 7104 27872
rect 7156 27860 7162 27872
rect 7300 27860 7328 28027
rect 9766 28024 9772 28027
rect 9824 28024 9830 28076
rect 11716 28074 12020 28094
rect 12051 28077 12109 28083
rect 12051 28074 12063 28077
rect 11716 28066 12063 28074
rect 11716 28064 11744 28066
rect 11440 28036 11744 28064
rect 11992 28046 12063 28066
rect 12051 28043 12063 28046
rect 12097 28043 12109 28077
rect 12051 28037 12109 28043
rect 8849 27999 8907 28005
rect 8849 27965 8861 27999
rect 8895 27996 8907 27999
rect 9030 27996 9036 28008
rect 8895 27968 9036 27996
rect 8895 27965 8907 27968
rect 8849 27959 8907 27965
rect 9030 27956 9036 27968
rect 9088 27956 9094 28008
rect 9398 27956 9404 28008
rect 9456 27996 9462 28008
rect 9585 27999 9643 28005
rect 9585 27996 9597 27999
rect 9456 27968 9597 27996
rect 9456 27956 9462 27968
rect 9585 27965 9597 27968
rect 9631 27965 9643 27999
rect 9585 27959 9643 27965
rect 9858 27956 9864 28008
rect 9916 27956 9922 28008
rect 8297 27931 8355 27937
rect 8297 27897 8309 27931
rect 8343 27928 8355 27931
rect 9309 27931 9367 27937
rect 9309 27928 9321 27931
rect 8343 27900 9321 27928
rect 8343 27897 8355 27900
rect 8297 27891 8355 27897
rect 9309 27897 9321 27900
rect 9355 27897 9367 27931
rect 9309 27891 9367 27897
rect 8110 27860 8116 27872
rect 7156 27832 8116 27860
rect 7156 27820 7162 27832
rect 8110 27820 8116 27832
rect 8168 27820 8174 27872
rect 8478 27820 8484 27872
rect 8536 27860 8542 27872
rect 9416 27860 9444 27956
rect 11054 27888 11060 27940
rect 11112 27928 11118 27940
rect 11440 27928 11468 28036
rect 12710 28024 12716 28076
rect 12768 28064 12774 28076
rect 13446 28073 13474 28104
rect 13814 28092 13820 28104
rect 13872 28092 13878 28144
rect 13173 28067 13231 28073
rect 13173 28064 13185 28067
rect 12768 28036 13185 28064
rect 12768 28024 12774 28036
rect 13173 28033 13185 28036
rect 13219 28033 13231 28067
rect 13173 28027 13231 28033
rect 13415 28067 13474 28073
rect 13415 28033 13427 28067
rect 13461 28036 13474 28067
rect 13461 28033 13473 28036
rect 13415 28027 13473 28033
rect 13538 28024 13544 28076
rect 13596 28064 13602 28076
rect 15562 28064 15568 28076
rect 13596 28036 15568 28064
rect 13596 28024 13602 28036
rect 15562 28024 15568 28036
rect 15620 28024 15626 28076
rect 11514 27956 11520 28008
rect 11572 27996 11578 28008
rect 11793 27999 11851 28005
rect 11793 27996 11805 27999
rect 11572 27968 11805 27996
rect 11572 27956 11578 27968
rect 11793 27965 11805 27968
rect 11839 27965 11851 27999
rect 11793 27959 11851 27965
rect 11606 27928 11612 27940
rect 11112 27900 11612 27928
rect 11112 27888 11118 27900
rect 11606 27888 11612 27900
rect 11664 27888 11670 27940
rect 12526 27860 12532 27872
rect 8536 27832 12532 27860
rect 8536 27820 8542 27832
rect 12526 27820 12532 27832
rect 12584 27820 12590 27872
rect 12802 27820 12808 27872
rect 12860 27820 12866 27872
rect 13170 27820 13176 27872
rect 13228 27860 13234 27872
rect 13538 27860 13544 27872
rect 13228 27832 13544 27860
rect 13228 27820 13234 27832
rect 13538 27820 13544 27832
rect 13596 27820 13602 27872
rect 13906 27820 13912 27872
rect 13964 27860 13970 27872
rect 14185 27863 14243 27869
rect 14185 27860 14197 27863
rect 13964 27832 14197 27860
rect 13964 27820 13970 27832
rect 14185 27829 14197 27832
rect 14231 27829 14243 27863
rect 14185 27823 14243 27829
rect 1104 27770 14812 27792
rect 1104 27718 2663 27770
rect 2715 27718 2727 27770
rect 2779 27718 2791 27770
rect 2843 27718 2855 27770
rect 2907 27718 2919 27770
rect 2971 27718 6090 27770
rect 6142 27718 6154 27770
rect 6206 27718 6218 27770
rect 6270 27718 6282 27770
rect 6334 27718 6346 27770
rect 6398 27718 9517 27770
rect 9569 27718 9581 27770
rect 9633 27718 9645 27770
rect 9697 27718 9709 27770
rect 9761 27718 9773 27770
rect 9825 27718 12944 27770
rect 12996 27718 13008 27770
rect 13060 27718 13072 27770
rect 13124 27718 13136 27770
rect 13188 27718 13200 27770
rect 13252 27718 14812 27770
rect 1104 27696 14812 27718
rect 7282 27656 7288 27668
rect 7024 27628 7288 27656
rect 5905 27591 5963 27597
rect 5905 27557 5917 27591
rect 5951 27588 5963 27591
rect 6917 27591 6975 27597
rect 6917 27588 6929 27591
rect 5951 27560 6929 27588
rect 5951 27557 5963 27560
rect 5905 27551 5963 27557
rect 6917 27557 6929 27560
rect 6963 27557 6975 27591
rect 6917 27551 6975 27557
rect 6457 27523 6515 27529
rect 6457 27489 6469 27523
rect 6503 27520 6515 27523
rect 6822 27520 6828 27532
rect 6503 27492 6828 27520
rect 6503 27489 6515 27492
rect 6457 27483 6515 27489
rect 6822 27480 6828 27492
rect 6880 27480 6886 27532
rect 7024 27520 7052 27628
rect 7282 27616 7288 27628
rect 7340 27616 7346 27668
rect 9858 27616 9864 27668
rect 9916 27656 9922 27668
rect 9953 27659 10011 27665
rect 9953 27656 9965 27659
rect 9916 27628 9965 27656
rect 9916 27616 9922 27628
rect 9953 27625 9965 27628
rect 9999 27625 10011 27659
rect 9953 27619 10011 27625
rect 12066 27616 12072 27668
rect 12124 27656 12130 27668
rect 15838 27656 15844 27668
rect 12124 27628 15844 27656
rect 12124 27616 12130 27628
rect 15838 27616 15844 27628
rect 15896 27616 15902 27668
rect 11606 27548 11612 27600
rect 11664 27588 11670 27600
rect 11664 27560 12204 27588
rect 11664 27548 11670 27560
rect 12176 27532 12204 27560
rect 13446 27548 13452 27600
rect 13504 27588 13510 27600
rect 13630 27588 13636 27600
rect 13504 27560 13636 27588
rect 13504 27548 13510 27560
rect 13630 27548 13636 27560
rect 13688 27548 13694 27600
rect 7193 27523 7251 27529
rect 7193 27520 7205 27523
rect 7024 27492 7205 27520
rect 7193 27489 7205 27492
rect 7239 27489 7251 27523
rect 7193 27483 7251 27489
rect 7310 27523 7368 27529
rect 7310 27489 7322 27523
rect 7356 27520 7368 27523
rect 7834 27520 7840 27532
rect 7356 27492 7840 27520
rect 7356 27489 7368 27492
rect 7310 27483 7368 27489
rect 7834 27480 7840 27492
rect 7892 27480 7898 27532
rect 8110 27480 8116 27532
rect 8168 27520 8174 27532
rect 8938 27520 8944 27532
rect 8168 27492 8944 27520
rect 8168 27480 8174 27492
rect 8938 27480 8944 27492
rect 8996 27480 9002 27532
rect 10134 27480 10140 27532
rect 10192 27520 10198 27532
rect 10318 27520 10324 27532
rect 10192 27492 10324 27520
rect 10192 27480 10198 27492
rect 10318 27480 10324 27492
rect 10376 27480 10382 27532
rect 11698 27480 11704 27532
rect 11756 27520 11762 27532
rect 11756 27492 12112 27520
rect 11756 27480 11762 27492
rect 4890 27412 4896 27464
rect 4948 27412 4954 27464
rect 6273 27455 6331 27461
rect 5151 27425 5209 27431
rect 750 27344 756 27396
rect 808 27384 814 27396
rect 1489 27387 1547 27393
rect 1489 27384 1501 27387
rect 808 27356 1501 27384
rect 808 27344 814 27356
rect 1489 27353 1501 27356
rect 1535 27353 1547 27387
rect 5151 27391 5163 27425
rect 5197 27422 5209 27425
rect 5197 27391 5212 27422
rect 6273 27421 6285 27455
rect 6319 27421 6331 27455
rect 6273 27415 6331 27421
rect 5151 27385 5212 27391
rect 5184 27384 5212 27385
rect 5258 27384 5264 27396
rect 5184 27356 5264 27384
rect 1489 27347 1547 27353
rect 5258 27344 5264 27356
rect 5316 27344 5322 27396
rect 1578 27276 1584 27328
rect 1636 27276 1642 27328
rect 6288 27316 6316 27415
rect 7466 27412 7472 27464
rect 7524 27412 7530 27464
rect 9214 27461 9220 27464
rect 9183 27455 9220 27461
rect 9183 27421 9195 27455
rect 9183 27415 9220 27421
rect 9214 27412 9220 27415
rect 9272 27412 9278 27464
rect 11977 27455 12035 27461
rect 11977 27452 11989 27455
rect 10060 27424 11989 27452
rect 8113 27387 8171 27393
rect 8113 27353 8125 27387
rect 8159 27384 8171 27387
rect 10060 27384 10088 27424
rect 11977 27421 11989 27424
rect 12023 27421 12035 27455
rect 12084 27452 12112 27492
rect 12158 27480 12164 27532
rect 12216 27480 12222 27532
rect 12434 27480 12440 27532
rect 12492 27520 12498 27532
rect 12621 27523 12679 27529
rect 12621 27520 12633 27523
rect 12492 27492 12633 27520
rect 12492 27480 12498 27492
rect 12621 27489 12633 27492
rect 12667 27489 12679 27523
rect 12621 27483 12679 27489
rect 12895 27455 12953 27461
rect 12895 27452 12907 27455
rect 12084 27424 12907 27452
rect 11977 27415 12035 27421
rect 12895 27421 12907 27424
rect 12941 27452 12953 27455
rect 13446 27452 13452 27464
rect 12941 27424 13452 27452
rect 12941 27421 12953 27424
rect 12895 27415 12953 27421
rect 13446 27412 13452 27424
rect 13504 27412 13510 27464
rect 8159 27356 10088 27384
rect 8159 27353 8171 27356
rect 8113 27347 8171 27353
rect 10134 27344 10140 27396
rect 10192 27384 10198 27396
rect 10873 27387 10931 27393
rect 10873 27384 10885 27387
rect 10192 27356 10885 27384
rect 10192 27344 10198 27356
rect 10873 27353 10885 27356
rect 10919 27353 10931 27387
rect 10873 27347 10931 27353
rect 11425 27387 11483 27393
rect 11425 27353 11437 27387
rect 11471 27384 11483 27387
rect 12345 27387 12403 27393
rect 11471 27356 11928 27384
rect 11471 27353 11483 27356
rect 11425 27347 11483 27353
rect 6730 27316 6736 27328
rect 6288 27288 6736 27316
rect 6730 27276 6736 27288
rect 6788 27276 6794 27328
rect 6822 27276 6828 27328
rect 6880 27316 6886 27328
rect 8202 27316 8208 27328
rect 6880 27288 8208 27316
rect 6880 27276 6886 27288
rect 8202 27276 8208 27288
rect 8260 27276 8266 27328
rect 11146 27276 11152 27328
rect 11204 27276 11210 27328
rect 11698 27276 11704 27328
rect 11756 27276 11762 27328
rect 11900 27316 11928 27356
rect 12345 27353 12357 27387
rect 12391 27384 12403 27387
rect 14182 27384 14188 27396
rect 12391 27356 14188 27384
rect 12391 27353 12403 27356
rect 12345 27347 12403 27353
rect 14182 27344 14188 27356
rect 14240 27344 14246 27396
rect 13262 27316 13268 27328
rect 11900 27288 13268 27316
rect 13262 27276 13268 27288
rect 13320 27276 13326 27328
rect 13633 27319 13691 27325
rect 13633 27285 13645 27319
rect 13679 27316 13691 27319
rect 13814 27316 13820 27328
rect 13679 27288 13820 27316
rect 13679 27285 13691 27288
rect 13633 27279 13691 27285
rect 13814 27276 13820 27288
rect 13872 27276 13878 27328
rect 1104 27226 14971 27248
rect 1104 27174 4376 27226
rect 4428 27174 4440 27226
rect 4492 27174 4504 27226
rect 4556 27174 4568 27226
rect 4620 27174 4632 27226
rect 4684 27174 7803 27226
rect 7855 27174 7867 27226
rect 7919 27174 7931 27226
rect 7983 27174 7995 27226
rect 8047 27174 8059 27226
rect 8111 27174 11230 27226
rect 11282 27174 11294 27226
rect 11346 27174 11358 27226
rect 11410 27174 11422 27226
rect 11474 27174 11486 27226
rect 11538 27174 14657 27226
rect 14709 27174 14721 27226
rect 14773 27174 14785 27226
rect 14837 27174 14849 27226
rect 14901 27174 14913 27226
rect 14965 27174 14971 27226
rect 1104 27152 14971 27174
rect 2961 27115 3019 27121
rect 2961 27081 2973 27115
rect 3007 27112 3019 27115
rect 3050 27112 3056 27124
rect 3007 27084 3056 27112
rect 3007 27081 3019 27084
rect 2961 27075 3019 27081
rect 3050 27072 3056 27084
rect 3108 27072 3114 27124
rect 5276 27084 8432 27112
rect 2777 26979 2835 26985
rect 2777 26945 2789 26979
rect 2823 26976 2835 26979
rect 3050 26976 3056 26988
rect 2823 26948 3056 26976
rect 2823 26945 2835 26948
rect 2777 26939 2835 26945
rect 3050 26936 3056 26948
rect 3108 26936 3114 26988
rect 4154 26936 4160 26988
rect 4212 26976 4218 26988
rect 5135 26979 5193 26985
rect 5135 26976 5147 26979
rect 4212 26948 5147 26976
rect 4212 26936 4218 26948
rect 5135 26945 5147 26948
rect 5181 26976 5193 26979
rect 5276 26976 5304 27084
rect 8404 27044 8432 27084
rect 8570 27072 8576 27124
rect 8628 27072 8634 27124
rect 8846 27072 8852 27124
rect 8904 27072 8910 27124
rect 11698 27072 11704 27124
rect 11756 27112 11762 27124
rect 14642 27112 14648 27124
rect 11756 27084 14648 27112
rect 11756 27072 11762 27084
rect 14642 27072 14648 27084
rect 14700 27072 14706 27124
rect 8864 27044 8892 27072
rect 8404 27016 8892 27044
rect 10686 27004 10692 27056
rect 10744 27004 10750 27056
rect 10962 27004 10968 27056
rect 11020 27044 11026 27056
rect 11020 27016 11744 27044
rect 11020 27004 11026 27016
rect 5181 26948 5304 26976
rect 5181 26945 5193 26948
rect 5135 26939 5193 26945
rect 5902 26936 5908 26988
rect 5960 26976 5966 26988
rect 6454 26976 6460 26988
rect 5960 26948 6460 26976
rect 5960 26936 5966 26948
rect 6454 26936 6460 26948
rect 6512 26936 6518 26988
rect 8570 26936 8576 26988
rect 8628 26976 8634 26988
rect 10195 26979 10253 26985
rect 10195 26976 10207 26979
rect 8628 26948 10207 26976
rect 8628 26936 8634 26948
rect 10195 26945 10207 26948
rect 10241 26945 10253 26979
rect 10704 26976 10732 27004
rect 11422 26976 11428 26988
rect 10704 26948 11428 26976
rect 10195 26939 10253 26945
rect 11422 26936 11428 26948
rect 11480 26976 11486 26988
rect 11517 26979 11575 26985
rect 11517 26976 11529 26979
rect 11480 26948 11529 26976
rect 11480 26936 11486 26948
rect 11517 26945 11529 26948
rect 11563 26945 11575 26979
rect 11517 26939 11575 26945
rect 11716 26920 11744 27016
rect 13354 27004 13360 27056
rect 13412 27004 13418 27056
rect 13722 27004 13728 27056
rect 13780 27004 13786 27056
rect 14090 27004 14096 27056
rect 14148 27004 14154 27056
rect 12434 26936 12440 26988
rect 12492 26936 12498 26988
rect 12710 26936 12716 26988
rect 12768 26936 12774 26988
rect 4890 26868 4896 26920
rect 4948 26868 4954 26920
rect 6730 26868 6736 26920
rect 6788 26868 6794 26920
rect 6822 26868 6828 26920
rect 6880 26908 6886 26920
rect 6917 26911 6975 26917
rect 6917 26908 6929 26911
rect 6880 26880 6929 26908
rect 6880 26868 6886 26880
rect 6917 26877 6929 26880
rect 6963 26877 6975 26911
rect 7653 26911 7711 26917
rect 7653 26908 7665 26911
rect 6917 26871 6975 26877
rect 7484 26880 7665 26908
rect 4908 26772 4936 26868
rect 5905 26843 5963 26849
rect 5905 26809 5917 26843
rect 5951 26840 5963 26843
rect 7377 26843 7435 26849
rect 7377 26840 7389 26843
rect 5951 26812 7389 26840
rect 5951 26809 5963 26812
rect 5905 26803 5963 26809
rect 7377 26809 7389 26812
rect 7423 26809 7435 26843
rect 7377 26803 7435 26809
rect 7098 26772 7104 26784
rect 4908 26744 7104 26772
rect 7098 26732 7104 26744
rect 7156 26732 7162 26784
rect 7484 26772 7512 26880
rect 7653 26877 7665 26880
rect 7699 26877 7711 26911
rect 7653 26871 7711 26877
rect 7742 26868 7748 26920
rect 7800 26917 7806 26920
rect 7800 26911 7828 26917
rect 7816 26877 7828 26911
rect 7800 26871 7828 26877
rect 7800 26868 7806 26871
rect 7926 26868 7932 26920
rect 7984 26868 7990 26920
rect 8938 26868 8944 26920
rect 8996 26908 9002 26920
rect 9858 26908 9864 26920
rect 8996 26880 9864 26908
rect 8996 26868 9002 26880
rect 9858 26868 9864 26880
rect 9916 26908 9922 26920
rect 9953 26911 10011 26917
rect 9953 26908 9965 26911
rect 9916 26880 9965 26908
rect 9916 26868 9922 26880
rect 9953 26877 9965 26880
rect 9999 26877 10011 26911
rect 9953 26871 10011 26877
rect 11698 26868 11704 26920
rect 11756 26868 11762 26920
rect 12575 26911 12633 26917
rect 12575 26877 12587 26911
rect 12621 26908 12633 26911
rect 12621 26880 13216 26908
rect 12621 26877 12633 26880
rect 12575 26871 12633 26877
rect 13188 26852 13216 26880
rect 9030 26800 9036 26852
rect 9088 26800 9094 26852
rect 10965 26843 11023 26849
rect 10965 26809 10977 26843
rect 11011 26840 11023 26843
rect 12161 26843 12219 26849
rect 12161 26840 12173 26843
rect 11011 26812 12173 26840
rect 11011 26809 11023 26812
rect 10965 26803 11023 26809
rect 12161 26809 12173 26812
rect 12207 26809 12219 26843
rect 12161 26803 12219 26809
rect 13170 26800 13176 26852
rect 13228 26840 13234 26852
rect 13354 26840 13360 26852
rect 13228 26812 13360 26840
rect 13228 26800 13234 26812
rect 13354 26800 13360 26812
rect 13412 26800 13418 26852
rect 9048 26772 9076 26800
rect 14108 26784 14136 27004
rect 7484 26744 9076 26772
rect 11514 26732 11520 26784
rect 11572 26772 11578 26784
rect 12710 26772 12716 26784
rect 11572 26744 12716 26772
rect 11572 26732 11578 26744
rect 12710 26732 12716 26744
rect 12768 26732 12774 26784
rect 13998 26732 14004 26784
rect 14056 26732 14062 26784
rect 14090 26732 14096 26784
rect 14148 26732 14154 26784
rect 1104 26682 14812 26704
rect 1104 26630 2663 26682
rect 2715 26630 2727 26682
rect 2779 26630 2791 26682
rect 2843 26630 2855 26682
rect 2907 26630 2919 26682
rect 2971 26630 6090 26682
rect 6142 26630 6154 26682
rect 6206 26630 6218 26682
rect 6270 26630 6282 26682
rect 6334 26630 6346 26682
rect 6398 26630 9517 26682
rect 9569 26630 9581 26682
rect 9633 26630 9645 26682
rect 9697 26630 9709 26682
rect 9761 26630 9773 26682
rect 9825 26630 12944 26682
rect 12996 26630 13008 26682
rect 13060 26630 13072 26682
rect 13124 26630 13136 26682
rect 13188 26630 13200 26682
rect 13252 26630 14812 26682
rect 1104 26608 14812 26630
rect 2869 26571 2927 26577
rect 2869 26537 2881 26571
rect 2915 26568 2927 26571
rect 3050 26568 3056 26580
rect 2915 26540 3056 26568
rect 2915 26537 2927 26540
rect 2869 26531 2927 26537
rect 3050 26528 3056 26540
rect 3108 26528 3114 26580
rect 7098 26568 7104 26580
rect 6748 26540 7104 26568
rect 1673 26503 1731 26509
rect 1673 26469 1685 26503
rect 1719 26500 1731 26503
rect 1719 26472 6666 26500
rect 1719 26469 1731 26472
rect 1673 26463 1731 26469
rect 3050 26324 3056 26376
rect 3108 26324 3114 26376
rect 6638 26364 6666 26472
rect 6748 26441 6776 26540
rect 7098 26528 7104 26540
rect 7156 26568 7162 26580
rect 7745 26571 7803 26577
rect 7156 26540 7512 26568
rect 7156 26528 7162 26540
rect 7484 26444 7512 26540
rect 7745 26537 7757 26571
rect 7791 26568 7803 26571
rect 7926 26568 7932 26580
rect 7791 26540 7932 26568
rect 7791 26537 7803 26540
rect 7745 26531 7803 26537
rect 7926 26528 7932 26540
rect 7984 26528 7990 26580
rect 10962 26528 10968 26580
rect 11020 26568 11026 26580
rect 11422 26568 11428 26580
rect 11020 26540 11428 26568
rect 11020 26528 11026 26540
rect 11422 26528 11428 26540
rect 11480 26528 11486 26580
rect 11514 26528 11520 26580
rect 11572 26528 11578 26580
rect 13262 26528 13268 26580
rect 13320 26568 13326 26580
rect 13909 26571 13967 26577
rect 13909 26568 13921 26571
rect 13320 26540 13921 26568
rect 13320 26528 13326 26540
rect 13909 26537 13921 26540
rect 13955 26537 13967 26571
rect 13909 26531 13967 26537
rect 12066 26460 12072 26512
rect 12124 26500 12130 26512
rect 12434 26500 12440 26512
rect 12124 26472 12440 26500
rect 12124 26460 12130 26472
rect 12434 26460 12440 26472
rect 12492 26460 12498 26512
rect 12713 26503 12771 26509
rect 12713 26469 12725 26503
rect 12759 26500 12771 26503
rect 12802 26500 12808 26512
rect 12759 26472 12808 26500
rect 12759 26469 12771 26472
rect 12713 26463 12771 26469
rect 12802 26460 12808 26472
rect 12860 26460 12866 26512
rect 6733 26435 6791 26441
rect 6733 26401 6745 26435
rect 6779 26401 6791 26435
rect 6733 26395 6791 26401
rect 7466 26392 7472 26444
rect 7524 26392 7530 26444
rect 9858 26392 9864 26444
rect 9916 26432 9922 26444
rect 9916 26404 10548 26432
rect 9916 26392 9922 26404
rect 6975 26367 7033 26373
rect 6975 26364 6987 26367
rect 6638 26336 6987 26364
rect 6975 26333 6987 26336
rect 7021 26364 7033 26367
rect 10226 26364 10232 26376
rect 7021 26336 10232 26364
rect 7021 26333 7033 26336
rect 6975 26327 7033 26333
rect 10226 26324 10232 26336
rect 10284 26324 10290 26376
rect 10520 26373 10548 26404
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 12989 26435 13047 26441
rect 12989 26432 13001 26435
rect 12676 26404 13001 26432
rect 12676 26392 12682 26404
rect 12989 26401 13001 26404
rect 13035 26401 13047 26435
rect 12989 26395 13047 26401
rect 13265 26435 13323 26441
rect 13265 26401 13277 26435
rect 13311 26432 13323 26435
rect 13906 26432 13912 26444
rect 13311 26404 13912 26432
rect 13311 26401 13323 26404
rect 13265 26395 13323 26401
rect 13906 26392 13912 26404
rect 13964 26392 13970 26444
rect 10505 26367 10563 26373
rect 10505 26333 10517 26367
rect 10551 26333 10563 26367
rect 10747 26367 10805 26373
rect 10747 26364 10759 26367
rect 10505 26327 10563 26333
rect 10612 26336 10759 26364
rect 1486 26256 1492 26308
rect 1544 26256 1550 26308
rect 1578 26256 1584 26308
rect 1636 26256 1642 26308
rect 8570 26296 8576 26308
rect 6746 26268 8576 26296
rect 1596 26228 1624 26256
rect 6746 26228 6774 26268
rect 8570 26256 8576 26268
rect 8628 26256 8634 26308
rect 8754 26256 8760 26308
rect 8812 26296 8818 26308
rect 10612 26296 10640 26336
rect 10747 26333 10759 26336
rect 10793 26333 10805 26367
rect 10747 26327 10805 26333
rect 12069 26367 12127 26373
rect 12069 26333 12081 26367
rect 12115 26364 12127 26367
rect 12158 26364 12164 26376
rect 12115 26336 12164 26364
rect 12115 26333 12127 26336
rect 12069 26327 12127 26333
rect 12158 26324 12164 26336
rect 12216 26324 12222 26376
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26364 12311 26367
rect 12434 26364 12440 26376
rect 12299 26336 12440 26364
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 12434 26324 12440 26336
rect 12492 26324 12498 26376
rect 13170 26373 13176 26376
rect 13127 26367 13176 26373
rect 13127 26333 13139 26367
rect 13173 26333 13176 26367
rect 13127 26327 13176 26333
rect 13170 26324 13176 26327
rect 13228 26324 13234 26376
rect 8812 26268 10640 26296
rect 8812 26256 8818 26268
rect 1596 26200 6774 26228
rect 15470 26188 15476 26240
rect 15528 26228 15534 26240
rect 15746 26228 15752 26240
rect 15528 26200 15752 26228
rect 15528 26188 15534 26200
rect 15746 26188 15752 26200
rect 15804 26188 15810 26240
rect 1104 26138 14971 26160
rect 1104 26086 4376 26138
rect 4428 26086 4440 26138
rect 4492 26086 4504 26138
rect 4556 26086 4568 26138
rect 4620 26086 4632 26138
rect 4684 26086 7803 26138
rect 7855 26086 7867 26138
rect 7919 26086 7931 26138
rect 7983 26086 7995 26138
rect 8047 26086 8059 26138
rect 8111 26086 11230 26138
rect 11282 26086 11294 26138
rect 11346 26086 11358 26138
rect 11410 26086 11422 26138
rect 11474 26086 11486 26138
rect 11538 26086 14657 26138
rect 14709 26086 14721 26138
rect 14773 26086 14785 26138
rect 14837 26086 14849 26138
rect 14901 26086 14913 26138
rect 14965 26086 14971 26138
rect 1104 26064 14971 26086
rect 13354 26024 13360 26036
rect 12176 25996 13360 26024
rect 5074 25916 5080 25968
rect 5132 25956 5138 25968
rect 12176 25965 12204 25996
rect 13354 25984 13360 25996
rect 13412 25984 13418 26036
rect 14090 25984 14096 26036
rect 14148 26024 14154 26036
rect 14461 26027 14519 26033
rect 14461 26024 14473 26027
rect 14148 25996 14473 26024
rect 14148 25984 14154 25996
rect 14461 25993 14473 25996
rect 14507 25993 14519 26027
rect 14461 25987 14519 25993
rect 12161 25959 12219 25965
rect 5132 25928 11652 25956
rect 5132 25916 5138 25928
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25888 1731 25891
rect 4154 25888 4160 25900
rect 1719 25860 4160 25888
rect 1719 25857 1731 25860
rect 1673 25851 1731 25857
rect 4154 25848 4160 25860
rect 4212 25848 4218 25900
rect 9859 25891 9917 25897
rect 9859 25857 9871 25891
rect 9905 25888 9917 25891
rect 10226 25888 10232 25900
rect 9905 25860 10232 25888
rect 9905 25857 9917 25860
rect 9859 25851 9917 25857
rect 10226 25848 10232 25860
rect 10284 25848 10290 25900
rect 11624 25897 11652 25928
rect 12161 25925 12173 25959
rect 12207 25925 12219 25959
rect 12161 25919 12219 25925
rect 11609 25891 11667 25897
rect 11609 25857 11621 25891
rect 11655 25857 11667 25891
rect 12805 25891 12863 25897
rect 12805 25888 12817 25891
rect 11609 25851 11667 25857
rect 12176 25860 12817 25888
rect 12176 25832 12204 25860
rect 12805 25857 12817 25860
rect 12851 25888 12863 25891
rect 12986 25888 12992 25900
rect 12851 25860 12992 25888
rect 12851 25857 12863 25860
rect 12805 25851 12863 25857
rect 12986 25848 12992 25860
rect 13044 25848 13050 25900
rect 13673 25897 13722 25898
rect 13673 25891 13737 25897
rect 13673 25857 13691 25891
rect 13725 25857 13737 25891
rect 13673 25851 13737 25857
rect 13673 25832 13701 25851
rect 13814 25848 13820 25900
rect 13872 25848 13878 25900
rect 750 25780 756 25832
rect 808 25820 814 25832
rect 1397 25823 1455 25829
rect 1397 25820 1409 25823
rect 808 25792 1409 25820
rect 808 25780 814 25792
rect 1397 25789 1409 25792
rect 1443 25789 1455 25823
rect 1397 25783 1455 25789
rect 9214 25780 9220 25832
rect 9272 25820 9278 25832
rect 9585 25823 9643 25829
rect 9585 25820 9597 25823
rect 9272 25792 9597 25820
rect 9272 25780 9278 25792
rect 9585 25789 9597 25792
rect 9631 25789 9643 25823
rect 9585 25783 9643 25789
rect 10686 25780 10692 25832
rect 10744 25820 10750 25832
rect 10962 25820 10968 25832
rect 10744 25792 10968 25820
rect 10744 25780 10750 25792
rect 10962 25780 10968 25792
rect 11020 25780 11026 25832
rect 12158 25780 12164 25832
rect 12216 25780 12222 25832
rect 12434 25780 12440 25832
rect 12492 25820 12498 25832
rect 12621 25823 12679 25829
rect 12621 25820 12633 25823
rect 12492 25792 12633 25820
rect 12492 25780 12498 25792
rect 12621 25789 12633 25792
rect 12667 25820 12679 25823
rect 12667 25792 12848 25820
rect 12667 25789 12679 25792
rect 12621 25783 12679 25789
rect 12820 25764 12848 25792
rect 13170 25780 13176 25832
rect 13228 25820 13234 25832
rect 13538 25820 13544 25832
rect 13228 25792 13544 25820
rect 13228 25780 13234 25792
rect 13538 25780 13544 25792
rect 13596 25780 13602 25832
rect 13630 25780 13636 25832
rect 13688 25792 13701 25832
rect 13688 25780 13694 25792
rect 12802 25712 12808 25764
rect 12860 25712 12866 25764
rect 13262 25712 13268 25764
rect 13320 25712 13326 25764
rect 10597 25687 10655 25693
rect 10597 25653 10609 25687
rect 10643 25684 10655 25687
rect 10962 25684 10968 25696
rect 10643 25656 10968 25684
rect 10643 25653 10655 25656
rect 10597 25647 10655 25653
rect 10962 25644 10968 25656
rect 11020 25644 11026 25696
rect 11882 25644 11888 25696
rect 11940 25644 11946 25696
rect 12437 25687 12495 25693
rect 12437 25653 12449 25687
rect 12483 25684 12495 25687
rect 14182 25684 14188 25696
rect 12483 25656 14188 25684
rect 12483 25653 12495 25656
rect 12437 25647 12495 25653
rect 14182 25644 14188 25656
rect 14240 25644 14246 25696
rect 1104 25594 14812 25616
rect 1104 25542 2663 25594
rect 2715 25542 2727 25594
rect 2779 25542 2791 25594
rect 2843 25542 2855 25594
rect 2907 25542 2919 25594
rect 2971 25542 6090 25594
rect 6142 25542 6154 25594
rect 6206 25542 6218 25594
rect 6270 25542 6282 25594
rect 6334 25542 6346 25594
rect 6398 25542 9517 25594
rect 9569 25542 9581 25594
rect 9633 25542 9645 25594
rect 9697 25542 9709 25594
rect 9761 25542 9773 25594
rect 9825 25542 12944 25594
rect 12996 25542 13008 25594
rect 13060 25542 13072 25594
rect 13124 25542 13136 25594
rect 13188 25542 13200 25594
rect 13252 25542 14812 25594
rect 1104 25520 14812 25542
rect 10594 25440 10600 25492
rect 10652 25440 10658 25492
rect 10778 25440 10784 25492
rect 10836 25440 10842 25492
rect 12342 25480 12348 25492
rect 11992 25452 12348 25480
rect 8481 25415 8539 25421
rect 8481 25381 8493 25415
rect 8527 25412 8539 25415
rect 9585 25415 9643 25421
rect 9585 25412 9597 25415
rect 8527 25384 9597 25412
rect 8527 25381 8539 25384
rect 8481 25375 8539 25381
rect 9585 25381 9597 25384
rect 9631 25381 9643 25415
rect 9585 25375 9643 25381
rect 9490 25304 9496 25356
rect 9548 25344 9554 25356
rect 10137 25347 10195 25353
rect 10137 25344 10149 25347
rect 9548 25316 10149 25344
rect 9548 25304 9554 25316
rect 10137 25313 10149 25316
rect 10183 25313 10195 25347
rect 10612 25344 10640 25440
rect 11992 25353 12020 25452
rect 12342 25440 12348 25452
rect 12400 25440 12406 25492
rect 12989 25483 13047 25489
rect 12989 25449 13001 25483
rect 13035 25480 13047 25483
rect 13262 25480 13268 25492
rect 13035 25452 13268 25480
rect 13035 25449 13047 25452
rect 12989 25443 13047 25449
rect 13262 25440 13268 25452
rect 13320 25440 13326 25492
rect 14550 25372 14556 25424
rect 14608 25412 14614 25424
rect 15562 25412 15568 25424
rect 14608 25384 15568 25412
rect 14608 25372 14614 25384
rect 15562 25372 15568 25384
rect 15620 25372 15626 25424
rect 11977 25347 12035 25353
rect 10612 25316 11192 25344
rect 10137 25307 10195 25313
rect 7098 25236 7104 25288
rect 7156 25236 7162 25288
rect 7374 25236 7380 25288
rect 7432 25276 7438 25288
rect 7469 25279 7527 25285
rect 7469 25276 7481 25279
rect 7432 25248 7481 25276
rect 7432 25236 7438 25248
rect 7469 25245 7481 25248
rect 7515 25245 7527 25279
rect 7469 25239 7527 25245
rect 7743 25279 7801 25285
rect 7743 25245 7755 25279
rect 7789 25276 7801 25279
rect 8202 25276 8208 25288
rect 7789 25248 8208 25276
rect 7789 25245 7801 25248
rect 7743 25239 7801 25245
rect 8202 25236 8208 25248
rect 8260 25236 8266 25288
rect 8478 25236 8484 25288
rect 8536 25276 8542 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8536 25248 8953 25276
rect 8536 25236 8542 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 7116 25208 7144 25236
rect 9140 25208 9168 25239
rect 9858 25236 9864 25288
rect 9916 25236 9922 25288
rect 9950 25236 9956 25288
rect 10008 25285 10014 25288
rect 10008 25279 10036 25285
rect 10024 25245 10036 25279
rect 11164 25276 11192 25316
rect 11977 25313 11989 25347
rect 12023 25313 12035 25347
rect 11977 25307 12035 25313
rect 12219 25279 12277 25285
rect 12219 25276 12231 25279
rect 11164 25248 12231 25276
rect 10008 25239 10036 25245
rect 12219 25245 12231 25248
rect 12265 25245 12277 25279
rect 12219 25239 12277 25245
rect 10008 25236 10014 25239
rect 11517 25211 11575 25217
rect 11517 25208 11529 25211
rect 7116 25180 9168 25208
rect 10612 25180 11529 25208
rect 8202 25100 8208 25152
rect 8260 25140 8266 25152
rect 10612 25140 10640 25180
rect 11517 25177 11529 25180
rect 11563 25177 11575 25211
rect 11517 25171 11575 25177
rect 11885 25211 11943 25217
rect 11885 25177 11897 25211
rect 11931 25208 11943 25211
rect 11974 25208 11980 25220
rect 11931 25180 11980 25208
rect 11931 25177 11943 25180
rect 11885 25171 11943 25177
rect 11974 25168 11980 25180
rect 12032 25168 12038 25220
rect 13538 25168 13544 25220
rect 13596 25168 13602 25220
rect 13906 25168 13912 25220
rect 13964 25168 13970 25220
rect 8260 25112 10640 25140
rect 8260 25100 8266 25112
rect 1104 25050 14971 25072
rect 1104 24998 4376 25050
rect 4428 24998 4440 25050
rect 4492 24998 4504 25050
rect 4556 24998 4568 25050
rect 4620 24998 4632 25050
rect 4684 24998 7803 25050
rect 7855 24998 7867 25050
rect 7919 24998 7931 25050
rect 7983 24998 7995 25050
rect 8047 24998 8059 25050
rect 8111 24998 11230 25050
rect 11282 24998 11294 25050
rect 11346 24998 11358 25050
rect 11410 24998 11422 25050
rect 11474 24998 11486 25050
rect 11538 24998 14657 25050
rect 14709 24998 14721 25050
rect 14773 24998 14785 25050
rect 14837 24998 14849 25050
rect 14901 24998 14913 25050
rect 14965 24998 14971 25050
rect 1104 24976 14971 24998
rect 7190 24896 7196 24948
rect 7248 24936 7254 24948
rect 7742 24936 7748 24948
rect 7248 24908 7748 24936
rect 7248 24896 7254 24908
rect 7742 24896 7748 24908
rect 7800 24896 7806 24948
rect 9490 24896 9496 24948
rect 9548 24896 9554 24948
rect 9858 24896 9864 24948
rect 9916 24936 9922 24948
rect 11238 24936 11244 24948
rect 9916 24908 11244 24936
rect 9916 24896 9922 24908
rect 11238 24896 11244 24908
rect 11296 24936 11302 24948
rect 12066 24936 12072 24948
rect 11296 24908 12072 24936
rect 11296 24896 11302 24908
rect 12066 24896 12072 24908
rect 12124 24896 12130 24948
rect 6546 24828 6552 24880
rect 6604 24828 6610 24880
rect 10244 24840 10548 24868
rect 750 24760 756 24812
rect 808 24800 814 24812
rect 1489 24803 1547 24809
rect 1489 24800 1501 24803
rect 808 24772 1501 24800
rect 808 24760 814 24772
rect 1489 24769 1501 24772
rect 1535 24769 1547 24803
rect 6564 24800 6592 24828
rect 1489 24763 1547 24769
rect 6472 24772 6592 24800
rect 5902 24692 5908 24744
rect 5960 24732 5966 24744
rect 6472 24741 6500 24772
rect 6638 24760 6644 24812
rect 6696 24800 6702 24812
rect 6731 24803 6789 24809
rect 6731 24800 6743 24803
rect 6696 24772 6743 24800
rect 6696 24760 6702 24772
rect 6731 24769 6743 24772
rect 6777 24769 6789 24803
rect 6731 24763 6789 24769
rect 7374 24760 7380 24812
rect 7432 24760 7438 24812
rect 7558 24760 7564 24812
rect 7616 24800 7622 24812
rect 8754 24809 8760 24812
rect 8723 24803 8760 24809
rect 8723 24800 8735 24803
rect 7616 24772 8735 24800
rect 7616 24760 7622 24772
rect 8723 24769 8735 24772
rect 8812 24800 8818 24812
rect 10244 24800 10272 24840
rect 8812 24772 10272 24800
rect 10319 24803 10377 24809
rect 8723 24763 8760 24769
rect 8754 24760 8760 24763
rect 8812 24760 8818 24772
rect 10319 24769 10331 24803
rect 10365 24800 10377 24803
rect 10410 24800 10416 24812
rect 10365 24772 10416 24800
rect 10365 24769 10377 24772
rect 10319 24763 10377 24769
rect 10410 24760 10416 24772
rect 10468 24760 10474 24812
rect 10520 24800 10548 24840
rect 11759 24803 11817 24809
rect 11759 24800 11771 24803
rect 10520 24772 11771 24800
rect 11759 24769 11771 24772
rect 11805 24769 11817 24803
rect 13170 24800 13176 24812
rect 13131 24772 13176 24800
rect 11759 24763 11817 24769
rect 13170 24760 13176 24772
rect 13228 24760 13234 24812
rect 6457 24735 6515 24741
rect 6457 24732 6469 24735
rect 5960 24704 6469 24732
rect 5960 24692 5966 24704
rect 6457 24701 6469 24704
rect 6503 24701 6515 24735
rect 7392 24732 7420 24760
rect 7926 24732 7932 24744
rect 7392 24704 7932 24732
rect 6457 24695 6515 24701
rect 7926 24692 7932 24704
rect 7984 24732 7990 24744
rect 8481 24735 8539 24741
rect 8481 24732 8493 24735
rect 7984 24704 8493 24732
rect 7984 24692 7990 24704
rect 8481 24701 8493 24704
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 9214 24692 9220 24744
rect 9272 24732 9278 24744
rect 10045 24735 10103 24741
rect 10045 24732 10057 24735
rect 9272 24704 10057 24732
rect 9272 24692 9278 24704
rect 10045 24701 10057 24704
rect 10091 24701 10103 24735
rect 11517 24735 11575 24741
rect 11517 24732 11529 24735
rect 10045 24695 10103 24701
rect 10704 24704 11529 24732
rect 1673 24667 1731 24673
rect 1673 24633 1685 24667
rect 1719 24664 1731 24667
rect 5534 24664 5540 24676
rect 1719 24636 5540 24664
rect 1719 24633 1731 24636
rect 1673 24627 1731 24633
rect 5534 24624 5540 24636
rect 5592 24624 5598 24676
rect 7374 24624 7380 24676
rect 7432 24664 7438 24676
rect 8386 24664 8392 24676
rect 7432 24636 8392 24664
rect 7432 24624 7438 24636
rect 8386 24624 8392 24636
rect 8444 24624 8450 24676
rect 7466 24556 7472 24608
rect 7524 24556 7530 24608
rect 7834 24556 7840 24608
rect 7892 24596 7898 24608
rect 8938 24596 8944 24608
rect 7892 24568 8944 24596
rect 7892 24556 7898 24568
rect 8938 24556 8944 24568
rect 8996 24596 9002 24608
rect 9858 24596 9864 24608
rect 8996 24568 9864 24596
rect 8996 24556 9002 24568
rect 9858 24556 9864 24568
rect 9916 24556 9922 24608
rect 10060 24596 10088 24695
rect 10704 24596 10732 24704
rect 11517 24701 11529 24704
rect 11563 24701 11575 24735
rect 12897 24735 12955 24741
rect 12897 24732 12909 24735
rect 11517 24695 11575 24701
rect 12406 24704 12909 24732
rect 11532 24608 11560 24695
rect 10060 24568 10732 24596
rect 11057 24599 11115 24605
rect 11057 24565 11069 24599
rect 11103 24596 11115 24599
rect 11422 24596 11428 24608
rect 11103 24568 11428 24596
rect 11103 24565 11115 24568
rect 11057 24559 11115 24565
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 11514 24556 11520 24608
rect 11572 24596 11578 24608
rect 12406 24596 12434 24704
rect 12897 24701 12909 24704
rect 12943 24701 12955 24735
rect 12897 24695 12955 24701
rect 11572 24568 12434 24596
rect 11572 24556 11578 24568
rect 12526 24556 12532 24608
rect 12584 24556 12590 24608
rect 13814 24556 13820 24608
rect 13872 24596 13878 24608
rect 13909 24599 13967 24605
rect 13909 24596 13921 24599
rect 13872 24568 13921 24596
rect 13872 24556 13878 24568
rect 13909 24565 13921 24568
rect 13955 24565 13967 24599
rect 13909 24559 13967 24565
rect 1104 24506 14812 24528
rect 1104 24454 2663 24506
rect 2715 24454 2727 24506
rect 2779 24454 2791 24506
rect 2843 24454 2855 24506
rect 2907 24454 2919 24506
rect 2971 24454 6090 24506
rect 6142 24454 6154 24506
rect 6206 24454 6218 24506
rect 6270 24454 6282 24506
rect 6334 24454 6346 24506
rect 6398 24454 9517 24506
rect 9569 24454 9581 24506
rect 9633 24454 9645 24506
rect 9697 24454 9709 24506
rect 9761 24454 9773 24506
rect 9825 24454 12944 24506
rect 12996 24454 13008 24506
rect 13060 24454 13072 24506
rect 13124 24454 13136 24506
rect 13188 24454 13200 24506
rect 13252 24454 14812 24506
rect 1104 24432 14812 24454
rect 7374 24392 7380 24404
rect 6288 24364 7380 24392
rect 4890 24148 4896 24200
rect 4948 24188 4954 24200
rect 5537 24191 5595 24197
rect 5537 24188 5549 24191
rect 4948 24160 5549 24188
rect 4948 24148 4954 24160
rect 5537 24157 5549 24160
rect 5583 24157 5595 24191
rect 5537 24151 5595 24157
rect 5811 24191 5869 24197
rect 5811 24157 5823 24191
rect 5857 24188 5869 24191
rect 6288 24188 6316 24364
rect 7374 24352 7380 24364
rect 7432 24352 7438 24404
rect 7466 24352 7472 24404
rect 7524 24392 7530 24404
rect 9953 24395 10011 24401
rect 9953 24392 9965 24395
rect 7524 24364 7604 24392
rect 7524 24352 7530 24364
rect 6730 24324 6736 24336
rect 6380 24296 6736 24324
rect 6380 24200 6408 24296
rect 6730 24284 6736 24296
rect 6788 24324 6794 24336
rect 7576 24333 7604 24364
rect 8588 24364 9965 24392
rect 7561 24327 7619 24333
rect 6788 24296 7328 24324
rect 6788 24284 6794 24296
rect 7300 24256 7328 24296
rect 7561 24293 7573 24327
rect 7607 24293 7619 24327
rect 7561 24287 7619 24293
rect 7954 24259 8012 24265
rect 7954 24256 7966 24259
rect 7300 24228 7966 24256
rect 7954 24225 7966 24228
rect 8000 24225 8012 24259
rect 7954 24219 8012 24225
rect 8113 24259 8171 24265
rect 8113 24225 8125 24259
rect 8159 24256 8171 24259
rect 8588 24256 8616 24364
rect 9953 24361 9965 24364
rect 9999 24361 10011 24395
rect 9953 24355 10011 24361
rect 11238 24352 11244 24404
rect 11296 24352 11302 24404
rect 11882 24352 11888 24404
rect 11940 24392 11946 24404
rect 12158 24392 12164 24404
rect 11940 24364 12164 24392
rect 11940 24352 11946 24364
rect 12158 24352 12164 24364
rect 12216 24352 12222 24404
rect 12526 24392 12532 24404
rect 12406 24364 12532 24392
rect 8159 24228 8616 24256
rect 8159 24225 8171 24228
rect 8113 24219 8171 24225
rect 8662 24216 8668 24268
rect 8720 24216 8726 24268
rect 11256 24256 11284 24352
rect 11422 24284 11428 24336
rect 11480 24284 11486 24336
rect 11882 24265 11888 24268
rect 11701 24259 11759 24265
rect 11701 24256 11713 24259
rect 11256 24228 11713 24256
rect 11701 24225 11713 24228
rect 11747 24225 11759 24259
rect 11701 24219 11759 24225
rect 11839 24259 11888 24265
rect 11839 24225 11851 24259
rect 11885 24225 11888 24259
rect 11839 24219 11888 24225
rect 11882 24216 11888 24219
rect 11940 24216 11946 24268
rect 11977 24259 12035 24265
rect 11977 24225 11989 24259
rect 12023 24256 12035 24259
rect 12406 24256 12434 24364
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 12621 24395 12679 24401
rect 12621 24361 12633 24395
rect 12667 24392 12679 24395
rect 13538 24392 13544 24404
rect 12667 24364 13544 24392
rect 12667 24361 12679 24364
rect 12621 24355 12679 24361
rect 13538 24352 13544 24364
rect 13596 24352 13602 24404
rect 12023 24228 12434 24256
rect 12023 24225 12035 24228
rect 11977 24219 12035 24225
rect 12618 24216 12624 24268
rect 12676 24256 12682 24268
rect 13538 24256 13544 24268
rect 12676 24228 13544 24256
rect 12676 24216 12682 24228
rect 13538 24216 13544 24228
rect 13596 24216 13602 24268
rect 5857 24160 6316 24188
rect 5857 24157 5869 24160
rect 5811 24151 5869 24157
rect 6362 24148 6368 24200
rect 6420 24148 6426 24200
rect 6730 24148 6736 24200
rect 6788 24188 6794 24200
rect 6917 24191 6975 24197
rect 6917 24188 6929 24191
rect 6788 24160 6929 24188
rect 6788 24148 6794 24160
rect 6917 24157 6929 24160
rect 6963 24157 6975 24191
rect 6917 24151 6975 24157
rect 7098 24148 7104 24200
rect 7156 24148 7162 24200
rect 7834 24148 7840 24200
rect 7892 24148 7898 24200
rect 8680 24188 8708 24216
rect 8941 24191 8999 24197
rect 8941 24188 8953 24191
rect 8680 24160 8953 24188
rect 8941 24157 8953 24160
rect 8987 24157 8999 24191
rect 8941 24151 8999 24157
rect 9122 24148 9128 24200
rect 9180 24188 9186 24200
rect 9215 24191 9273 24197
rect 9215 24188 9227 24191
rect 9180 24160 9227 24188
rect 9180 24148 9186 24160
rect 9215 24157 9227 24160
rect 9261 24157 9273 24191
rect 9215 24151 9273 24157
rect 9306 24148 9312 24200
rect 9364 24148 9370 24200
rect 10778 24148 10784 24200
rect 10836 24148 10842 24200
rect 10965 24191 11023 24197
rect 10965 24157 10977 24191
rect 11011 24157 11023 24191
rect 10965 24151 11023 24157
rect 750 24080 756 24132
rect 808 24120 814 24132
rect 1489 24123 1547 24129
rect 1489 24120 1501 24123
rect 808 24092 1501 24120
rect 808 24080 814 24092
rect 1489 24089 1501 24092
rect 1535 24089 1547 24123
rect 1489 24083 1547 24089
rect 1673 24123 1731 24129
rect 1673 24089 1685 24123
rect 1719 24120 1731 24123
rect 4982 24120 4988 24132
rect 1719 24092 4988 24120
rect 1719 24089 1731 24092
rect 1673 24083 1731 24089
rect 4982 24080 4988 24092
rect 5040 24080 5046 24132
rect 8662 24080 8668 24132
rect 8720 24120 8726 24132
rect 9140 24120 9168 24148
rect 8720 24092 9168 24120
rect 8720 24080 8726 24092
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 7558 24052 7564 24064
rect 6595 24024 7564 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 8757 24055 8815 24061
rect 8757 24021 8769 24055
rect 8803 24052 8815 24055
rect 9324 24052 9352 24148
rect 8803 24024 9352 24052
rect 10980 24052 11008 24151
rect 13170 24080 13176 24132
rect 13228 24080 13234 24132
rect 13541 24123 13599 24129
rect 13541 24089 13553 24123
rect 13587 24120 13599 24123
rect 15102 24120 15108 24132
rect 13587 24092 15108 24120
rect 13587 24089 13599 24092
rect 13541 24083 13599 24089
rect 15102 24080 15108 24092
rect 15160 24080 15166 24132
rect 11698 24052 11704 24064
rect 10980 24024 11704 24052
rect 8803 24021 8815 24024
rect 8757 24015 8815 24021
rect 11698 24012 11704 24024
rect 11756 24052 11762 24064
rect 13262 24052 13268 24064
rect 11756 24024 13268 24052
rect 11756 24012 11762 24024
rect 13262 24012 13268 24024
rect 13320 24012 13326 24064
rect 13354 24012 13360 24064
rect 13412 24052 13418 24064
rect 13722 24052 13728 24064
rect 13412 24024 13728 24052
rect 13412 24012 13418 24024
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 1104 23962 14971 23984
rect 1104 23910 4376 23962
rect 4428 23910 4440 23962
rect 4492 23910 4504 23962
rect 4556 23910 4568 23962
rect 4620 23910 4632 23962
rect 4684 23910 7803 23962
rect 7855 23910 7867 23962
rect 7919 23910 7931 23962
rect 7983 23910 7995 23962
rect 8047 23910 8059 23962
rect 8111 23910 11230 23962
rect 11282 23910 11294 23962
rect 11346 23910 11358 23962
rect 11410 23910 11422 23962
rect 11474 23910 11486 23962
rect 11538 23910 14657 23962
rect 14709 23910 14721 23962
rect 14773 23910 14785 23962
rect 14837 23910 14849 23962
rect 14901 23910 14913 23962
rect 14965 23910 14971 23962
rect 1104 23888 14971 23910
rect 6822 23848 6828 23860
rect 6564 23820 6828 23848
rect 3050 23672 3056 23724
rect 3108 23712 3114 23724
rect 4890 23712 4896 23724
rect 3108 23684 4896 23712
rect 3108 23672 3114 23684
rect 4890 23672 4896 23684
rect 4948 23672 4954 23724
rect 5166 23712 5172 23724
rect 5127 23684 5172 23712
rect 5166 23672 5172 23684
rect 5224 23672 5230 23724
rect 6564 23721 6592 23820
rect 6822 23808 6828 23820
rect 6880 23848 6886 23860
rect 6880 23820 8064 23848
rect 6880 23808 6886 23820
rect 8036 23780 8064 23820
rect 8202 23808 8208 23860
rect 8260 23808 8266 23860
rect 13170 23808 13176 23860
rect 13228 23848 13234 23860
rect 13228 23820 14320 23848
rect 13228 23808 13234 23820
rect 10226 23780 10232 23792
rect 8036 23752 10232 23780
rect 10226 23740 10232 23752
rect 10284 23740 10290 23792
rect 10778 23740 10784 23792
rect 10836 23780 10842 23792
rect 12526 23780 12532 23792
rect 10836 23752 12532 23780
rect 10836 23740 10842 23752
rect 12526 23740 12532 23752
rect 12584 23740 12590 23792
rect 14292 23780 14320 23820
rect 14461 23783 14519 23789
rect 14461 23780 14473 23783
rect 14292 23752 14473 23780
rect 14461 23749 14473 23752
rect 14507 23749 14519 23783
rect 14461 23743 14519 23749
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 7282 23672 7288 23724
rect 7340 23672 7346 23724
rect 7558 23672 7564 23724
rect 7616 23672 7622 23724
rect 8846 23672 8852 23724
rect 8904 23712 8910 23724
rect 9367 23715 9425 23721
rect 9367 23712 9379 23715
rect 8904 23684 9379 23712
rect 8904 23672 8910 23684
rect 9367 23681 9379 23684
rect 9413 23681 9425 23715
rect 9367 23675 9425 23681
rect 12158 23672 12164 23724
rect 12216 23672 12222 23724
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23681 12679 23715
rect 12621 23675 12679 23681
rect 4908 23508 4936 23672
rect 5994 23604 6000 23656
rect 6052 23644 6058 23656
rect 6362 23644 6368 23656
rect 6052 23616 6368 23644
rect 6052 23604 6058 23616
rect 6362 23604 6368 23616
rect 6420 23604 6426 23656
rect 7374 23604 7380 23656
rect 7432 23653 7438 23656
rect 7432 23647 7460 23653
rect 7448 23613 7460 23647
rect 7432 23607 7460 23613
rect 9125 23647 9183 23653
rect 9125 23613 9137 23647
rect 9171 23613 9183 23647
rect 9125 23607 9183 23613
rect 7432 23604 7438 23607
rect 5905 23579 5963 23585
rect 5905 23545 5917 23579
rect 5951 23576 5963 23579
rect 7009 23579 7067 23585
rect 7009 23576 7021 23579
rect 5951 23548 7021 23576
rect 5951 23545 5963 23548
rect 5905 23539 5963 23545
rect 7009 23545 7021 23548
rect 7055 23545 7067 23579
rect 7009 23539 7067 23545
rect 9140 23508 9168 23607
rect 12066 23604 12072 23656
rect 12124 23644 12130 23656
rect 12250 23644 12256 23656
rect 12124 23616 12256 23644
rect 12124 23604 12130 23616
rect 12250 23604 12256 23616
rect 12308 23644 12314 23656
rect 12634 23644 12662 23675
rect 13814 23672 13820 23724
rect 13872 23672 13878 23724
rect 12308 23616 12662 23644
rect 12308 23604 12314 23616
rect 12802 23604 12808 23656
rect 12860 23604 12866 23656
rect 13538 23604 13544 23656
rect 13596 23604 13602 23656
rect 13630 23604 13636 23656
rect 13688 23653 13694 23656
rect 13688 23647 13716 23653
rect 13704 23613 13716 23647
rect 13688 23607 13716 23613
rect 13688 23604 13694 23607
rect 13262 23536 13268 23588
rect 13320 23536 13326 23588
rect 9214 23508 9220 23520
rect 4908 23480 9220 23508
rect 9214 23468 9220 23480
rect 9272 23468 9278 23520
rect 10134 23468 10140 23520
rect 10192 23468 10198 23520
rect 12437 23511 12495 23517
rect 12437 23477 12449 23511
rect 12483 23508 12495 23511
rect 14182 23508 14188 23520
rect 12483 23480 14188 23508
rect 12483 23477 12495 23480
rect 12437 23471 12495 23477
rect 14182 23468 14188 23480
rect 14240 23468 14246 23520
rect 1104 23418 14812 23440
rect 1104 23366 2663 23418
rect 2715 23366 2727 23418
rect 2779 23366 2791 23418
rect 2843 23366 2855 23418
rect 2907 23366 2919 23418
rect 2971 23366 6090 23418
rect 6142 23366 6154 23418
rect 6206 23366 6218 23418
rect 6270 23366 6282 23418
rect 6334 23366 6346 23418
rect 6398 23366 9517 23418
rect 9569 23366 9581 23418
rect 9633 23366 9645 23418
rect 9697 23366 9709 23418
rect 9761 23366 9773 23418
rect 9825 23366 12944 23418
rect 12996 23366 13008 23418
rect 13060 23366 13072 23418
rect 13124 23366 13136 23418
rect 13188 23366 13200 23418
rect 13252 23366 14812 23418
rect 1104 23344 14812 23366
rect 5442 23264 5448 23316
rect 5500 23304 5506 23316
rect 7190 23304 7196 23316
rect 5500 23276 7196 23304
rect 5500 23264 5506 23276
rect 7190 23264 7196 23276
rect 7248 23264 7254 23316
rect 7282 23264 7288 23316
rect 7340 23304 7346 23316
rect 7466 23304 7472 23316
rect 7340 23276 7472 23304
rect 7340 23264 7346 23276
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 11977 23307 12035 23313
rect 11977 23273 11989 23307
rect 12023 23304 12035 23307
rect 12710 23304 12716 23316
rect 12023 23276 12716 23304
rect 12023 23273 12035 23276
rect 11977 23267 12035 23273
rect 12710 23264 12716 23276
rect 12768 23264 12774 23316
rect 13262 23264 13268 23316
rect 13320 23304 13326 23316
rect 13357 23307 13415 23313
rect 13357 23304 13369 23307
rect 13320 23276 13369 23304
rect 13320 23264 13326 23276
rect 13357 23273 13369 23276
rect 13403 23273 13415 23307
rect 13357 23267 13415 23273
rect 9398 23128 9404 23180
rect 9456 23168 9462 23180
rect 10965 23171 11023 23177
rect 10965 23168 10977 23171
rect 9456 23140 10977 23168
rect 9456 23128 9462 23140
rect 10965 23137 10977 23140
rect 11011 23137 11023 23171
rect 10965 23131 11023 23137
rect 11698 23128 11704 23180
rect 11756 23168 11762 23180
rect 11974 23168 11980 23180
rect 11756 23140 11980 23168
rect 11756 23128 11762 23140
rect 11974 23128 11980 23140
rect 12032 23168 12038 23180
rect 12345 23171 12403 23177
rect 12345 23168 12357 23171
rect 12032 23140 12357 23168
rect 12032 23128 12038 23140
rect 12345 23137 12357 23140
rect 12391 23137 12403 23171
rect 12345 23131 12403 23137
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 8846 23100 8852 23112
rect 1719 23072 8852 23100
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 8846 23060 8852 23072
rect 8904 23060 8910 23112
rect 10870 23060 10876 23112
rect 10928 23060 10934 23112
rect 11146 23060 11152 23112
rect 11204 23100 11210 23112
rect 11239 23103 11297 23109
rect 11239 23100 11251 23103
rect 11204 23072 11251 23100
rect 11204 23060 11210 23072
rect 11239 23069 11251 23072
rect 11285 23069 11297 23103
rect 12618 23100 12624 23112
rect 12579 23072 12624 23100
rect 11239 23063 11297 23069
rect 12618 23060 12624 23072
rect 12676 23060 12682 23112
rect 14185 23103 14243 23109
rect 14185 23069 14197 23103
rect 14231 23100 14243 23103
rect 14366 23100 14372 23112
rect 14231 23072 14372 23100
rect 14231 23069 14243 23072
rect 14185 23063 14243 23069
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 750 22992 756 23044
rect 808 23032 814 23044
rect 1489 23035 1547 23041
rect 1489 23032 1501 23035
rect 808 23004 1501 23032
rect 808 22992 814 23004
rect 1489 23001 1501 23004
rect 1535 23001 1547 23035
rect 10888 23032 10916 23060
rect 12986 23032 12992 23044
rect 10888 23004 12992 23032
rect 1489 22995 1547 23001
rect 12986 22992 12992 23004
rect 13044 22992 13050 23044
rect 10502 22924 10508 22976
rect 10560 22964 10566 22976
rect 12618 22964 12624 22976
rect 10560 22936 12624 22964
rect 10560 22924 10566 22936
rect 12618 22924 12624 22936
rect 12676 22964 12682 22976
rect 12802 22964 12808 22976
rect 12676 22936 12808 22964
rect 12676 22924 12682 22936
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 14369 22967 14427 22973
rect 14369 22933 14381 22967
rect 14415 22964 14427 22967
rect 15102 22964 15108 22976
rect 14415 22936 15108 22964
rect 14415 22933 14427 22936
rect 14369 22927 14427 22933
rect 15102 22924 15108 22936
rect 15160 22924 15166 22976
rect 15286 22896 15292 22908
rect 1104 22874 14971 22896
rect 1104 22822 4376 22874
rect 4428 22822 4440 22874
rect 4492 22822 4504 22874
rect 4556 22822 4568 22874
rect 4620 22822 4632 22874
rect 4684 22822 7803 22874
rect 7855 22822 7867 22874
rect 7919 22822 7931 22874
rect 7983 22822 7995 22874
rect 8047 22822 8059 22874
rect 8111 22822 11230 22874
rect 11282 22822 11294 22874
rect 11346 22822 11358 22874
rect 11410 22822 11422 22874
rect 11474 22822 11486 22874
rect 11538 22822 14657 22874
rect 14709 22822 14721 22874
rect 14773 22822 14785 22874
rect 14837 22822 14849 22874
rect 14901 22822 14913 22874
rect 14965 22822 14971 22874
rect 1104 22800 14971 22822
rect 15028 22868 15292 22896
rect 1581 22763 1639 22769
rect 1581 22729 1593 22763
rect 1627 22760 1639 22763
rect 1670 22760 1676 22772
rect 1627 22732 1676 22760
rect 1627 22729 1639 22732
rect 1581 22723 1639 22729
rect 1670 22720 1676 22732
rect 1728 22760 1734 22772
rect 2314 22760 2320 22772
rect 1728 22732 2320 22760
rect 1728 22720 1734 22732
rect 2314 22720 2320 22732
rect 2372 22720 2378 22772
rect 10318 22720 10324 22772
rect 10376 22720 10382 22772
rect 12986 22720 12992 22772
rect 13044 22760 13050 22772
rect 13357 22763 13415 22769
rect 13357 22760 13369 22763
rect 13044 22732 13369 22760
rect 13044 22720 13050 22732
rect 13357 22729 13369 22732
rect 13403 22729 13415 22763
rect 13538 22760 13544 22772
rect 13357 22723 13415 22729
rect 13464 22732 13544 22760
rect 10336 22692 10364 22720
rect 10334 22664 10364 22692
rect 10334 22663 10362 22664
rect 10303 22657 10362 22663
rect 750 22584 756 22636
rect 808 22624 814 22636
rect 1489 22627 1547 22633
rect 1489 22624 1501 22627
rect 808 22596 1501 22624
rect 808 22584 814 22596
rect 1489 22593 1501 22596
rect 1535 22593 1547 22627
rect 8386 22624 8392 22636
rect 8347 22596 8392 22624
rect 1489 22587 1547 22593
rect 8386 22584 8392 22596
rect 8444 22584 8450 22636
rect 9398 22584 9404 22636
rect 9456 22624 9462 22636
rect 10045 22627 10103 22633
rect 10045 22624 10057 22627
rect 9456 22596 10057 22624
rect 9456 22584 9462 22596
rect 10045 22593 10057 22596
rect 10091 22593 10103 22627
rect 10303 22623 10315 22657
rect 10349 22626 10362 22657
rect 12618 22633 12624 22636
rect 11701 22627 11759 22633
rect 10349 22623 10361 22626
rect 11701 22624 11713 22627
rect 10303 22617 10361 22623
rect 10045 22587 10103 22593
rect 10796 22596 11713 22624
rect 10796 22568 10824 22596
rect 11701 22593 11713 22596
rect 11747 22593 11759 22627
rect 12437 22627 12495 22633
rect 12437 22624 12449 22627
rect 11701 22587 11759 22593
rect 12434 22593 12449 22624
rect 12483 22593 12495 22627
rect 12434 22587 12495 22593
rect 12575 22627 12624 22633
rect 12575 22593 12587 22627
rect 12621 22593 12624 22627
rect 12575 22587 12624 22593
rect 7742 22516 7748 22568
rect 7800 22556 7806 22568
rect 8113 22559 8171 22565
rect 8113 22556 8125 22559
rect 7800 22528 8125 22556
rect 7800 22516 7806 22528
rect 8113 22525 8125 22528
rect 8159 22525 8171 22559
rect 8113 22519 8171 22525
rect 10778 22516 10784 22568
rect 10836 22516 10842 22568
rect 10870 22516 10876 22568
rect 10928 22556 10934 22568
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 10928 22528 11529 22556
rect 10928 22516 10934 22528
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 12434 22556 12462 22587
rect 12618 22584 12624 22587
rect 12676 22584 12682 22636
rect 12710 22584 12716 22636
rect 12768 22584 12774 22636
rect 11517 22519 11575 22525
rect 12268 22528 12462 22556
rect 11057 22491 11115 22497
rect 11057 22457 11069 22491
rect 11103 22488 11115 22491
rect 12161 22491 12219 22497
rect 12161 22488 12173 22491
rect 11103 22460 12173 22488
rect 11103 22457 11115 22460
rect 11057 22451 11115 22457
rect 12161 22457 12173 22460
rect 12207 22457 12219 22491
rect 12161 22451 12219 22457
rect 9122 22380 9128 22432
rect 9180 22380 9186 22432
rect 9398 22380 9404 22432
rect 9456 22420 9462 22432
rect 12268 22420 12296 22528
rect 13464 22420 13492 22732
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 14274 22720 14280 22772
rect 14332 22760 14338 22772
rect 14369 22763 14427 22769
rect 14369 22760 14381 22763
rect 14332 22732 14381 22760
rect 14332 22720 14338 22732
rect 14369 22729 14381 22732
rect 14415 22729 14427 22763
rect 14369 22723 14427 22729
rect 14918 22720 14924 22772
rect 14976 22760 14982 22772
rect 15028 22760 15056 22868
rect 15286 22856 15292 22868
rect 15344 22856 15350 22908
rect 15102 22788 15108 22840
rect 15160 22828 15166 22840
rect 15470 22828 15476 22840
rect 15160 22800 15476 22828
rect 15160 22788 15166 22800
rect 15470 22788 15476 22800
rect 15528 22788 15534 22840
rect 14976 22732 15056 22760
rect 14976 22720 14982 22732
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 15252 22732 15424 22760
rect 15252 22720 15258 22732
rect 15396 22704 15424 22732
rect 15378 22652 15384 22704
rect 15436 22652 15442 22704
rect 13538 22584 13544 22636
rect 13596 22584 13602 22636
rect 14093 22627 14151 22633
rect 14093 22593 14105 22627
rect 14139 22624 14151 22627
rect 15930 22624 15936 22636
rect 14139 22596 15936 22624
rect 14139 22593 14151 22596
rect 14093 22587 14151 22593
rect 15930 22584 15936 22596
rect 15988 22584 15994 22636
rect 13722 22516 13728 22568
rect 13780 22556 13786 22568
rect 15654 22556 15660 22568
rect 13780 22528 15660 22556
rect 13780 22516 13786 22528
rect 15654 22516 15660 22528
rect 15712 22516 15718 22568
rect 14918 22448 14924 22500
rect 14976 22488 14982 22500
rect 15286 22488 15292 22500
rect 14976 22460 15292 22488
rect 14976 22448 14982 22460
rect 15286 22448 15292 22460
rect 15344 22448 15350 22500
rect 9456 22392 13492 22420
rect 9456 22380 9462 22392
rect 13814 22380 13820 22432
rect 13872 22380 13878 22432
rect 14366 22380 14372 22432
rect 14424 22420 14430 22432
rect 15562 22420 15568 22432
rect 14424 22392 15568 22420
rect 14424 22380 14430 22392
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 1104 22330 14812 22352
rect 1104 22278 2663 22330
rect 2715 22278 2727 22330
rect 2779 22278 2791 22330
rect 2843 22278 2855 22330
rect 2907 22278 2919 22330
rect 2971 22278 6090 22330
rect 6142 22278 6154 22330
rect 6206 22278 6218 22330
rect 6270 22278 6282 22330
rect 6334 22278 6346 22330
rect 6398 22278 9517 22330
rect 9569 22278 9581 22330
rect 9633 22278 9645 22330
rect 9697 22278 9709 22330
rect 9761 22278 9773 22330
rect 9825 22278 12944 22330
rect 12996 22278 13008 22330
rect 13060 22278 13072 22330
rect 13124 22278 13136 22330
rect 13188 22278 13200 22330
rect 13252 22278 14812 22330
rect 1104 22256 14812 22278
rect 5166 22176 5172 22228
rect 5224 22216 5230 22228
rect 7742 22216 7748 22228
rect 5224 22188 6684 22216
rect 5224 22176 5230 22188
rect 5534 21972 5540 22024
rect 5592 21972 5598 22024
rect 5902 21972 5908 22024
rect 5960 22012 5966 22024
rect 6270 22021 6276 22024
rect 5997 22015 6055 22021
rect 5997 22012 6009 22015
rect 5960 21984 6009 22012
rect 5960 21972 5966 21984
rect 5997 21981 6009 21984
rect 6043 21981 6055 22015
rect 6239 22015 6276 22021
rect 6239 22012 6251 22015
rect 5997 21975 6055 21981
rect 6086 21984 6251 22012
rect 5552 21944 5580 21972
rect 6086 21944 6114 21984
rect 6239 21981 6251 21984
rect 6239 21975 6276 21981
rect 6270 21972 6276 21975
rect 6328 21972 6334 22024
rect 6656 22012 6684 22188
rect 7392 22188 7748 22216
rect 7392 22089 7420 22188
rect 7742 22176 7748 22188
rect 7800 22176 7806 22228
rect 10778 22216 10784 22228
rect 9784 22188 10784 22216
rect 9030 22108 9036 22160
rect 9088 22148 9094 22160
rect 9088 22120 9674 22148
rect 9088 22108 9094 22120
rect 7377 22083 7435 22089
rect 7377 22049 7389 22083
rect 7423 22049 7435 22083
rect 7377 22043 7435 22049
rect 7558 22012 7564 22024
rect 6656 21984 7564 22012
rect 7558 21972 7564 21984
rect 7616 22012 7622 22024
rect 7651 22015 7709 22021
rect 7651 22012 7663 22015
rect 7616 21984 7663 22012
rect 7616 21972 7622 21984
rect 7651 21981 7663 21984
rect 7697 21981 7709 22015
rect 9646 22012 9674 22120
rect 9784 22092 9812 22188
rect 10778 22176 10784 22188
rect 10836 22176 10842 22228
rect 11882 22176 11888 22228
rect 11940 22216 11946 22228
rect 12894 22216 12900 22228
rect 11940 22188 12900 22216
rect 11940 22176 11946 22188
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 13446 22176 13452 22228
rect 13504 22216 13510 22228
rect 13630 22216 13636 22228
rect 13504 22188 13636 22216
rect 13504 22176 13510 22188
rect 13630 22176 13636 22188
rect 13688 22176 13694 22228
rect 14274 22176 14280 22228
rect 14332 22176 14338 22228
rect 10318 22148 10324 22160
rect 9874 22120 10324 22148
rect 9766 22040 9772 22092
rect 9824 22040 9830 22092
rect 9874 22012 9902 22120
rect 10318 22108 10324 22120
rect 10376 22108 10382 22160
rect 10134 22040 10140 22092
rect 10192 22080 10198 22092
rect 10413 22083 10471 22089
rect 10413 22080 10425 22083
rect 10192 22052 10425 22080
rect 10192 22040 10198 22052
rect 10413 22049 10425 22052
rect 10459 22049 10471 22083
rect 10413 22043 10471 22049
rect 10502 22040 10508 22092
rect 10560 22080 10566 22092
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 10560 22052 10701 22080
rect 10560 22040 10566 22052
rect 10689 22049 10701 22052
rect 10735 22049 10747 22083
rect 10689 22043 10747 22049
rect 10962 22040 10968 22092
rect 11020 22040 11026 22092
rect 10870 22021 10876 22024
rect 9646 21984 9902 22012
rect 9953 22015 10011 22021
rect 7651 21975 7709 21981
rect 9953 21981 9965 22015
rect 9999 21981 10011 22015
rect 9953 21975 10011 21981
rect 10827 22015 10876 22021
rect 10827 21981 10839 22015
rect 10873 21981 10876 22015
rect 10827 21975 10876 21981
rect 5552 21916 6114 21944
rect 7009 21879 7067 21885
rect 7009 21845 7021 21879
rect 7055 21876 7067 21879
rect 7558 21876 7564 21888
rect 7055 21848 7564 21876
rect 7055 21845 7067 21848
rect 7009 21839 7067 21845
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 8386 21836 8392 21888
rect 8444 21836 8450 21888
rect 9968 21876 9996 21975
rect 10870 21972 10876 21975
rect 10928 21972 10934 22024
rect 11974 21972 11980 22024
rect 12032 22012 12038 22024
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 12032 21984 12173 22012
rect 12032 21972 12038 21984
rect 12161 21981 12173 21984
rect 12207 21981 12219 22015
rect 12419 21985 12477 21991
rect 12419 21982 12431 21985
rect 12161 21975 12219 21981
rect 12406 21951 12431 21982
rect 12465 21951 12477 21985
rect 12894 21972 12900 22024
rect 12952 22012 12958 22024
rect 14093 22015 14151 22021
rect 12952 21984 14044 22012
rect 12952 21972 12958 21984
rect 12406 21945 12477 21951
rect 12406 21944 12434 21945
rect 13446 21944 13452 21956
rect 11532 21916 12434 21944
rect 12728 21916 13452 21944
rect 10318 21876 10324 21888
rect 9968 21848 10324 21876
rect 10318 21836 10324 21848
rect 10376 21836 10382 21888
rect 10686 21836 10692 21888
rect 10744 21876 10750 21888
rect 11532 21876 11560 21916
rect 10744 21848 11560 21876
rect 10744 21836 10750 21848
rect 11606 21836 11612 21888
rect 11664 21836 11670 21888
rect 12434 21836 12440 21888
rect 12492 21876 12498 21888
rect 12728 21876 12756 21916
rect 13446 21904 13452 21916
rect 13504 21904 13510 21956
rect 14016 21944 14044 21984
rect 14093 21981 14105 22015
rect 14139 22012 14151 22015
rect 14274 22012 14280 22024
rect 14139 21984 14280 22012
rect 14139 21981 14151 21984
rect 14093 21975 14151 21981
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 15838 21944 15844 21956
rect 14016 21916 15844 21944
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 12492 21848 12756 21876
rect 13173 21879 13231 21885
rect 12492 21836 12498 21848
rect 13173 21845 13185 21879
rect 13219 21876 13231 21879
rect 13262 21876 13268 21888
rect 13219 21848 13268 21876
rect 13219 21845 13231 21848
rect 13173 21839 13231 21845
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 1104 21786 14971 21808
rect 1104 21734 4376 21786
rect 4428 21734 4440 21786
rect 4492 21734 4504 21786
rect 4556 21734 4568 21786
rect 4620 21734 4632 21786
rect 4684 21734 7803 21786
rect 7855 21734 7867 21786
rect 7919 21734 7931 21786
rect 7983 21734 7995 21786
rect 8047 21734 8059 21786
rect 8111 21734 11230 21786
rect 11282 21734 11294 21786
rect 11346 21734 11358 21786
rect 11410 21734 11422 21786
rect 11474 21734 11486 21786
rect 11538 21734 14657 21786
rect 14709 21734 14721 21786
rect 14773 21734 14785 21786
rect 14837 21734 14849 21786
rect 14901 21734 14913 21786
rect 14965 21734 14971 21786
rect 1104 21712 14971 21734
rect 4982 21632 4988 21684
rect 5040 21672 5046 21684
rect 5040 21644 9812 21672
rect 5040 21632 5046 21644
rect 6656 21575 6684 21644
rect 6623 21569 6684 21575
rect 750 21496 756 21548
rect 808 21536 814 21548
rect 1489 21539 1547 21545
rect 1489 21536 1501 21539
rect 808 21508 1501 21536
rect 808 21496 814 21508
rect 1489 21505 1501 21508
rect 1535 21505 1547 21539
rect 6623 21535 6635 21569
rect 6669 21538 6684 21569
rect 6822 21564 6828 21616
rect 6880 21604 6886 21616
rect 7098 21604 7104 21616
rect 6880 21576 7104 21604
rect 6880 21564 6886 21576
rect 7098 21564 7104 21576
rect 7156 21564 7162 21616
rect 7466 21564 7472 21616
rect 7524 21604 7530 21616
rect 7926 21604 7932 21616
rect 7524 21576 7932 21604
rect 7524 21564 7530 21576
rect 7926 21564 7932 21576
rect 7984 21564 7990 21616
rect 9784 21604 9812 21644
rect 9858 21632 9864 21684
rect 9916 21632 9922 21684
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12434 21672 12440 21684
rect 11931 21644 12440 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12434 21632 12440 21644
rect 12492 21632 12498 21684
rect 13722 21672 13728 21684
rect 12544 21644 13728 21672
rect 10686 21604 10692 21616
rect 9784 21576 10692 21604
rect 10686 21564 10692 21576
rect 10744 21564 10750 21616
rect 12544 21613 12572 21644
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 12529 21607 12587 21613
rect 12529 21573 12541 21607
rect 12575 21573 12587 21607
rect 12529 21567 12587 21573
rect 8205 21539 8263 21545
rect 6669 21535 6681 21538
rect 8205 21536 8217 21539
rect 6623 21529 6681 21535
rect 1489 21499 1547 21505
rect 7852 21508 8217 21536
rect 7852 21480 7880 21508
rect 8205 21505 8217 21508
rect 8251 21505 8263 21539
rect 8205 21502 8263 21505
rect 8205 21499 8294 21502
rect 5902 21428 5908 21480
rect 5960 21468 5966 21480
rect 6365 21471 6423 21477
rect 6365 21468 6377 21471
rect 5960 21440 6377 21468
rect 5960 21428 5966 21440
rect 6365 21437 6377 21440
rect 6411 21437 6423 21471
rect 6365 21431 6423 21437
rect 7834 21428 7840 21480
rect 7892 21428 7898 21480
rect 8018 21428 8024 21480
rect 8076 21428 8082 21480
rect 8220 21474 8294 21499
rect 8386 21496 8392 21548
rect 8444 21496 8450 21548
rect 9214 21496 9220 21548
rect 9272 21496 9278 21548
rect 10870 21496 10876 21548
rect 10928 21536 10934 21548
rect 11609 21539 11667 21545
rect 11609 21536 11621 21539
rect 10928 21508 11621 21536
rect 10928 21496 10934 21508
rect 11609 21505 11621 21508
rect 11655 21505 11667 21539
rect 11609 21499 11667 21505
rect 12158 21496 12164 21548
rect 12216 21496 12222 21548
rect 13541 21539 13599 21545
rect 12268 21508 13032 21536
rect 8266 21468 8294 21474
rect 8404 21468 8432 21496
rect 12268 21480 12296 21508
rect 8665 21471 8723 21477
rect 8665 21468 8677 21471
rect 8266 21440 8340 21468
rect 8404 21440 8677 21468
rect 1673 21403 1731 21409
rect 1673 21369 1685 21403
rect 1719 21369 1731 21403
rect 1673 21363 1731 21369
rect 7300 21372 7512 21400
rect 1688 21332 1716 21363
rect 7300 21332 7328 21372
rect 1688 21304 7328 21332
rect 7374 21292 7380 21344
rect 7432 21292 7438 21344
rect 7484 21332 7512 21372
rect 8202 21332 8208 21344
rect 7484 21304 8208 21332
rect 8202 21292 8208 21304
rect 8260 21292 8266 21344
rect 8312 21332 8340 21440
rect 8665 21437 8677 21440
rect 8711 21437 8723 21471
rect 8665 21431 8723 21437
rect 8754 21428 8760 21480
rect 8812 21468 8818 21480
rect 8938 21468 8944 21480
rect 8812 21440 8944 21468
rect 8812 21428 8818 21440
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 9122 21477 9128 21480
rect 9079 21471 9128 21477
rect 9079 21437 9091 21471
rect 9125 21437 9128 21471
rect 9079 21431 9128 21437
rect 9122 21428 9128 21431
rect 9180 21468 9186 21480
rect 12250 21468 12256 21480
rect 9180 21440 12256 21468
rect 9180 21428 9186 21440
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 12621 21471 12679 21477
rect 12621 21468 12633 21471
rect 12406 21440 12633 21468
rect 12406 21400 12434 21440
rect 12621 21437 12633 21440
rect 12667 21437 12679 21471
rect 12621 21431 12679 21437
rect 12805 21471 12863 21477
rect 12805 21437 12817 21471
rect 12851 21468 12863 21471
rect 12894 21468 12900 21480
rect 12851 21440 12900 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 9968 21372 12434 21400
rect 13004 21400 13032 21508
rect 13541 21505 13553 21539
rect 13587 21505 13599 21539
rect 13541 21499 13599 21505
rect 13262 21428 13268 21480
rect 13320 21428 13326 21480
rect 13556 21468 13584 21499
rect 13372 21440 13584 21468
rect 13372 21400 13400 21440
rect 13630 21428 13636 21480
rect 13688 21477 13694 21480
rect 13688 21471 13716 21477
rect 13704 21437 13716 21471
rect 13688 21431 13716 21437
rect 13688 21428 13694 21431
rect 13814 21428 13820 21480
rect 13872 21428 13878 21480
rect 14458 21428 14464 21480
rect 14516 21468 14522 21480
rect 15930 21468 15936 21480
rect 14516 21440 15936 21468
rect 14516 21428 14522 21440
rect 15930 21428 15936 21440
rect 15988 21428 15994 21480
rect 13004 21372 13400 21400
rect 9968 21332 9996 21372
rect 8312 21304 9996 21332
rect 10686 21292 10692 21344
rect 10744 21332 10750 21344
rect 10962 21332 10968 21344
rect 10744 21304 10968 21332
rect 10744 21292 10750 21304
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 14274 21332 14280 21344
rect 12492 21304 14280 21332
rect 12492 21292 12498 21304
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14461 21335 14519 21341
rect 14461 21301 14473 21335
rect 14507 21332 14519 21335
rect 14507 21304 14872 21332
rect 14507 21301 14519 21304
rect 14461 21295 14519 21301
rect 1104 21242 14812 21264
rect 1104 21190 2663 21242
rect 2715 21190 2727 21242
rect 2779 21190 2791 21242
rect 2843 21190 2855 21242
rect 2907 21190 2919 21242
rect 2971 21190 6090 21242
rect 6142 21190 6154 21242
rect 6206 21190 6218 21242
rect 6270 21190 6282 21242
rect 6334 21190 6346 21242
rect 6398 21190 9517 21242
rect 9569 21190 9581 21242
rect 9633 21190 9645 21242
rect 9697 21190 9709 21242
rect 9761 21190 9773 21242
rect 9825 21190 12944 21242
rect 12996 21190 13008 21242
rect 13060 21190 13072 21242
rect 13124 21190 13136 21242
rect 13188 21190 13200 21242
rect 13252 21190 14812 21242
rect 1104 21168 14812 21190
rect 3326 21088 3332 21140
rect 3384 21088 3390 21140
rect 7374 21128 7380 21140
rect 7116 21100 7380 21128
rect 3234 21020 3240 21072
rect 3292 21060 3298 21072
rect 6546 21060 6552 21072
rect 3292 21032 6552 21060
rect 3292 21020 3298 21032
rect 6546 21020 6552 21032
rect 6604 21060 6610 21072
rect 6730 21060 6736 21072
rect 6604 21032 6736 21060
rect 6604 21020 6610 21032
rect 6730 21020 6736 21032
rect 6788 21020 6794 21072
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20992 1731 20995
rect 6914 20992 6920 21004
rect 1719 20964 6920 20992
rect 1719 20961 1731 20964
rect 1673 20955 1731 20961
rect 6914 20952 6920 20964
rect 6972 20952 6978 21004
rect 7009 20995 7067 21001
rect 7009 20961 7021 20995
rect 7055 20992 7067 20995
rect 7116 20992 7144 21100
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 7650 21088 7656 21140
rect 7708 21128 7714 21140
rect 8205 21131 8263 21137
rect 8205 21128 8217 21131
rect 7708 21100 8217 21128
rect 7708 21088 7714 21100
rect 8205 21097 8217 21100
rect 8251 21097 8263 21131
rect 11885 21131 11943 21137
rect 8205 21091 8263 21097
rect 9876 21100 11560 21128
rect 8018 21020 8024 21072
rect 8076 21060 8082 21072
rect 9876 21060 9904 21100
rect 8076 21032 9904 21060
rect 8076 21020 8082 21032
rect 7055 20964 7144 20992
rect 7285 20995 7343 21001
rect 7055 20961 7067 20964
rect 7009 20955 7067 20961
rect 7285 20961 7297 20995
rect 7331 20992 7343 20995
rect 7926 20992 7932 21004
rect 7331 20964 7932 20992
rect 7331 20961 7343 20964
rect 7285 20955 7343 20961
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 2498 20884 2504 20936
rect 2556 20924 2562 20936
rect 3145 20927 3203 20933
rect 3145 20924 3157 20927
rect 2556 20896 3157 20924
rect 2556 20884 2562 20896
rect 3145 20893 3157 20896
rect 3191 20893 3203 20927
rect 3145 20887 3203 20893
rect 6365 20927 6423 20933
rect 6365 20893 6377 20927
rect 6411 20924 6423 20927
rect 6454 20924 6460 20936
rect 6411 20896 6460 20924
rect 6411 20893 6423 20896
rect 6365 20887 6423 20893
rect 6454 20884 6460 20896
rect 6512 20884 6518 20936
rect 6546 20884 6552 20936
rect 6604 20884 6610 20936
rect 7374 20884 7380 20936
rect 7432 20933 7438 20936
rect 7432 20927 7460 20933
rect 7448 20893 7460 20927
rect 7432 20887 7460 20893
rect 7432 20884 7438 20887
rect 7558 20884 7564 20936
rect 7616 20884 7622 20936
rect 8266 20868 8294 21032
rect 8570 20884 8576 20936
rect 8628 20884 8634 20936
rect 9766 20884 9772 20936
rect 9824 20884 9830 20936
rect 10011 20927 10069 20933
rect 10011 20924 10023 20927
rect 9993 20893 10023 20924
rect 10057 20893 10069 20927
rect 9993 20887 10069 20893
rect 8202 20816 8208 20868
rect 8260 20828 8294 20868
rect 8588 20856 8616 20884
rect 9674 20856 9680 20868
rect 8588 20828 9680 20856
rect 8260 20816 8266 20828
rect 9674 20816 9680 20828
rect 9732 20816 9738 20868
rect 6730 20748 6736 20800
rect 6788 20788 6794 20800
rect 9993 20788 10021 20887
rect 10502 20884 10508 20936
rect 10560 20924 10566 20936
rect 11425 20927 11483 20933
rect 11425 20924 11437 20927
rect 10560 20896 11437 20924
rect 10560 20884 10566 20896
rect 11425 20893 11437 20896
rect 11471 20893 11483 20927
rect 11425 20887 11483 20893
rect 6788 20760 10021 20788
rect 6788 20748 6794 20760
rect 10778 20748 10784 20800
rect 10836 20748 10842 20800
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 11241 20791 11299 20797
rect 11241 20788 11253 20791
rect 11204 20760 11253 20788
rect 11204 20748 11210 20760
rect 11241 20757 11253 20760
rect 11287 20757 11299 20791
rect 11532 20788 11560 21100
rect 11885 21097 11897 21131
rect 11931 21128 11943 21131
rect 13633 21131 13691 21137
rect 11931 21100 13584 21128
rect 11931 21097 11943 21100
rect 11885 21091 11943 21097
rect 13556 21060 13584 21100
rect 13633 21097 13645 21131
rect 13679 21128 13691 21131
rect 13814 21128 13820 21140
rect 13679 21100 13820 21128
rect 13679 21097 13691 21100
rect 13633 21091 13691 21097
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 14090 21060 14096 21072
rect 13556 21032 14096 21060
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 11974 20952 11980 21004
rect 12032 20992 12038 21004
rect 12250 20992 12256 21004
rect 12032 20964 12256 20992
rect 12032 20952 12038 20964
rect 12250 20952 12256 20964
rect 12308 20992 12314 21004
rect 12621 20995 12679 21001
rect 12621 20992 12633 20995
rect 12308 20964 12633 20992
rect 12308 20952 12314 20964
rect 12621 20961 12633 20964
rect 12667 20961 12679 20995
rect 12621 20955 12679 20961
rect 12894 20933 12900 20936
rect 11609 20927 11667 20933
rect 11609 20893 11621 20927
rect 11655 20924 11667 20927
rect 12879 20927 12900 20933
rect 11655 20896 12848 20924
rect 11655 20893 11667 20896
rect 11609 20887 11667 20893
rect 12158 20816 12164 20868
rect 12216 20816 12222 20868
rect 12526 20816 12532 20868
rect 12584 20816 12590 20868
rect 12820 20856 12848 20896
rect 12879 20893 12891 20927
rect 12879 20887 12900 20893
rect 12894 20884 12900 20887
rect 12952 20884 12958 20936
rect 14844 20856 14872 21304
rect 12820 20828 14872 20856
rect 13630 20788 13636 20800
rect 11532 20760 13636 20788
rect 11241 20751 11299 20757
rect 13630 20748 13636 20760
rect 13688 20788 13694 20800
rect 13688 20760 15976 20788
rect 13688 20748 13694 20760
rect 15948 20732 15976 20760
rect 1104 20698 14971 20720
rect 1104 20646 4376 20698
rect 4428 20646 4440 20698
rect 4492 20646 4504 20698
rect 4556 20646 4568 20698
rect 4620 20646 4632 20698
rect 4684 20646 7803 20698
rect 7855 20646 7867 20698
rect 7919 20646 7931 20698
rect 7983 20646 7995 20698
rect 8047 20646 8059 20698
rect 8111 20646 11230 20698
rect 11282 20646 11294 20698
rect 11346 20646 11358 20698
rect 11410 20646 11422 20698
rect 11474 20646 11486 20698
rect 11538 20646 14657 20698
rect 14709 20646 14721 20698
rect 14773 20646 14785 20698
rect 14837 20646 14849 20698
rect 14901 20646 14913 20698
rect 14965 20646 14971 20698
rect 15930 20680 15936 20732
rect 15988 20680 15994 20732
rect 1104 20624 14971 20646
rect 4982 20544 4988 20596
rect 5040 20544 5046 20596
rect 7009 20587 7067 20593
rect 7009 20553 7021 20587
rect 7055 20553 7067 20587
rect 7009 20547 7067 20553
rect 5000 20448 5028 20544
rect 7024 20516 7052 20547
rect 7926 20544 7932 20596
rect 7984 20584 7990 20596
rect 7984 20556 10732 20584
rect 7984 20544 7990 20556
rect 9398 20516 9404 20528
rect 7024 20488 7512 20516
rect 5057 20451 5115 20457
rect 5057 20448 5069 20451
rect 5000 20420 5069 20448
rect 5057 20417 5069 20420
rect 5103 20448 5115 20451
rect 6457 20451 6515 20457
rect 6457 20448 6469 20451
rect 5103 20420 6469 20448
rect 5103 20417 5115 20420
rect 5057 20411 5115 20417
rect 6457 20417 6469 20420
rect 6503 20417 6515 20451
rect 6457 20411 6515 20417
rect 7193 20451 7251 20457
rect 7193 20417 7205 20451
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 4798 20340 4804 20392
rect 4856 20340 4862 20392
rect 6641 20383 6699 20389
rect 6641 20349 6653 20383
rect 6687 20380 6699 20383
rect 7208 20380 7236 20411
rect 7282 20408 7288 20460
rect 7340 20408 7346 20460
rect 7484 20457 7512 20488
rect 7576 20488 9404 20516
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20417 7527 20451
rect 7469 20411 7527 20417
rect 7576 20380 7604 20488
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 9674 20476 9680 20528
rect 9732 20516 9738 20528
rect 10502 20516 10508 20528
rect 9732 20488 10508 20516
rect 9732 20476 9738 20488
rect 10502 20476 10508 20488
rect 10560 20476 10566 20528
rect 8386 20408 8392 20460
rect 8444 20448 8450 20460
rect 8479 20451 8537 20457
rect 8479 20448 8491 20451
rect 8444 20420 8491 20448
rect 8444 20408 8450 20420
rect 8479 20417 8491 20420
rect 8525 20448 8537 20451
rect 9827 20451 9885 20457
rect 9827 20448 9839 20451
rect 8525 20420 9839 20448
rect 8525 20417 8537 20420
rect 8479 20411 8537 20417
rect 9827 20417 9839 20420
rect 9873 20417 9885 20451
rect 9827 20411 9885 20417
rect 6687 20352 7604 20380
rect 6687 20349 6699 20352
rect 6641 20343 6699 20349
rect 7926 20340 7932 20392
rect 7984 20380 7990 20392
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 7984 20352 8217 20380
rect 7984 20340 7990 20352
rect 8205 20349 8217 20352
rect 8251 20349 8263 20383
rect 8205 20343 8263 20349
rect 9398 20340 9404 20392
rect 9456 20380 9462 20392
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 9456 20352 9597 20380
rect 9456 20340 9462 20352
rect 9585 20349 9597 20352
rect 9631 20349 9643 20383
rect 10704 20380 10732 20556
rect 11146 20544 11152 20596
rect 11204 20544 11210 20596
rect 11977 20587 12035 20593
rect 11977 20553 11989 20587
rect 12023 20584 12035 20587
rect 13906 20584 13912 20596
rect 12023 20556 13912 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 14001 20587 14059 20593
rect 14001 20553 14013 20587
rect 14047 20584 14059 20587
rect 15194 20584 15200 20596
rect 14047 20556 15200 20584
rect 14047 20553 14059 20556
rect 14001 20547 14059 20553
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 10778 20476 10784 20528
rect 10836 20476 10842 20528
rect 11164 20516 11192 20544
rect 11164 20488 11376 20516
rect 10796 20448 10824 20476
rect 11146 20448 11152 20460
rect 10796 20420 11152 20448
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 11348 20457 11376 20488
rect 11606 20476 11612 20528
rect 11664 20516 11670 20528
rect 13725 20519 13783 20525
rect 13725 20516 13737 20519
rect 11664 20488 13737 20516
rect 11664 20476 11670 20488
rect 13725 20485 13737 20488
rect 13771 20485 13783 20519
rect 13725 20479 13783 20485
rect 11333 20451 11391 20457
rect 11333 20417 11345 20451
rect 11379 20417 11391 20451
rect 11333 20411 11391 20417
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 10704 20352 11560 20380
rect 9585 20343 9643 20349
rect 6181 20315 6239 20321
rect 6181 20281 6193 20315
rect 6227 20312 6239 20315
rect 11330 20312 11336 20324
rect 6227 20284 8340 20312
rect 6227 20281 6239 20284
rect 6181 20275 6239 20281
rect 7006 20204 7012 20256
rect 7064 20244 7070 20256
rect 7190 20244 7196 20256
rect 7064 20216 7196 20244
rect 7064 20204 7070 20216
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 7374 20204 7380 20256
rect 7432 20204 7438 20256
rect 8312 20244 8340 20284
rect 10520 20284 11336 20312
rect 8570 20244 8576 20256
rect 8312 20216 8576 20244
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 9214 20204 9220 20256
rect 9272 20204 9278 20256
rect 9306 20204 9312 20256
rect 9364 20244 9370 20256
rect 10520 20244 10548 20284
rect 11330 20272 11336 20284
rect 11388 20272 11394 20324
rect 11532 20312 11560 20352
rect 11606 20340 11612 20392
rect 11664 20380 11670 20392
rect 11716 20380 11744 20411
rect 12342 20408 12348 20460
rect 12400 20448 12406 20460
rect 12435 20451 12493 20457
rect 12435 20448 12447 20451
rect 12400 20420 12447 20448
rect 12400 20408 12406 20420
rect 12435 20417 12447 20420
rect 12481 20417 12493 20451
rect 12435 20411 12493 20417
rect 11664 20352 11744 20380
rect 12161 20383 12219 20389
rect 11664 20340 11670 20352
rect 12161 20349 12173 20383
rect 12207 20349 12219 20383
rect 12161 20343 12219 20349
rect 12176 20312 12204 20343
rect 11532 20284 12204 20312
rect 9364 20216 10548 20244
rect 10597 20247 10655 20253
rect 9364 20204 9370 20216
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 11054 20244 11060 20256
rect 10643 20216 11060 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11241 20247 11299 20253
rect 11241 20213 11253 20247
rect 11287 20244 11299 20247
rect 11698 20244 11704 20256
rect 11287 20216 11704 20244
rect 11287 20213 11299 20216
rect 11241 20207 11299 20213
rect 11698 20204 11704 20216
rect 11756 20204 11762 20256
rect 12176 20244 12204 20284
rect 12250 20244 12256 20256
rect 12176 20216 12256 20244
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 12618 20204 12624 20256
rect 12676 20244 12682 20256
rect 13173 20247 13231 20253
rect 13173 20244 13185 20247
rect 12676 20216 13185 20244
rect 12676 20204 12682 20216
rect 13173 20213 13185 20216
rect 13219 20213 13231 20247
rect 13173 20207 13231 20213
rect 1104 20154 14812 20176
rect 1104 20102 2663 20154
rect 2715 20102 2727 20154
rect 2779 20102 2791 20154
rect 2843 20102 2855 20154
rect 2907 20102 2919 20154
rect 2971 20102 6090 20154
rect 6142 20102 6154 20154
rect 6206 20102 6218 20154
rect 6270 20102 6282 20154
rect 6334 20102 6346 20154
rect 6398 20102 9517 20154
rect 9569 20102 9581 20154
rect 9633 20102 9645 20154
rect 9697 20102 9709 20154
rect 9761 20102 9773 20154
rect 9825 20102 12944 20154
rect 12996 20102 13008 20154
rect 13060 20102 13072 20154
rect 13124 20102 13136 20154
rect 13188 20102 13200 20154
rect 13252 20102 14812 20154
rect 1104 20080 14812 20102
rect 2406 20000 2412 20052
rect 2464 20040 2470 20052
rect 7926 20040 7932 20052
rect 2464 20012 7420 20040
rect 2464 20000 2470 20012
rect 1673 19975 1731 19981
rect 1673 19941 1685 19975
rect 1719 19972 1731 19975
rect 5534 19972 5540 19984
rect 1719 19944 5540 19972
rect 1719 19941 1731 19944
rect 1673 19935 1731 19941
rect 5534 19932 5540 19944
rect 5592 19932 5598 19984
rect 5810 19932 5816 19984
rect 5868 19932 5874 19984
rect 6825 19975 6883 19981
rect 6825 19941 6837 19975
rect 6871 19972 6883 19975
rect 7282 19972 7288 19984
rect 6871 19944 7288 19972
rect 6871 19941 6883 19944
rect 6825 19935 6883 19941
rect 5828 19904 5856 19932
rect 5736 19876 5856 19904
rect 750 19728 756 19780
rect 808 19768 814 19780
rect 1489 19771 1547 19777
rect 1489 19768 1501 19771
rect 808 19740 1501 19768
rect 808 19728 814 19740
rect 1489 19737 1501 19740
rect 1535 19737 1547 19771
rect 1489 19731 1547 19737
rect 1118 19660 1124 19712
rect 1176 19700 1182 19712
rect 5736 19700 5764 19876
rect 7116 19848 7144 19944
rect 7282 19932 7288 19944
rect 7340 19932 7346 19984
rect 5810 19796 5816 19848
rect 5868 19796 5874 19848
rect 6087 19829 6145 19835
rect 6087 19795 6099 19829
rect 6133 19795 6145 19829
rect 6914 19796 6920 19848
rect 6972 19796 6978 19848
rect 7098 19796 7104 19848
rect 7156 19796 7162 19848
rect 7392 19845 7420 20012
rect 7484 20012 7932 20040
rect 7484 19913 7512 20012
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 9214 20000 9220 20052
rect 9272 20040 9278 20052
rect 10781 20043 10839 20049
rect 9272 20012 10548 20040
rect 9272 20000 9278 20012
rect 8481 19975 8539 19981
rect 8481 19941 8493 19975
rect 8527 19972 8539 19975
rect 9585 19975 9643 19981
rect 9585 19972 9597 19975
rect 8527 19944 9597 19972
rect 8527 19941 8539 19944
rect 8481 19935 8539 19941
rect 9585 19941 9597 19944
rect 9631 19941 9643 19975
rect 9585 19935 9643 19941
rect 7469 19907 7527 19913
rect 7469 19873 7481 19907
rect 7515 19873 7527 19907
rect 7469 19867 7527 19873
rect 8938 19864 8944 19916
rect 8996 19864 9002 19916
rect 9856 19864 9862 19916
rect 9914 19904 9920 19916
rect 10135 19907 10193 19913
rect 9914 19876 9959 19904
rect 9914 19864 9920 19876
rect 10135 19873 10147 19907
rect 10181 19904 10193 19907
rect 10520 19904 10548 20012
rect 10781 20009 10793 20043
rect 10827 20040 10839 20043
rect 10870 20040 10876 20052
rect 10827 20012 10876 20040
rect 10827 20009 10839 20012
rect 10781 20003 10839 20009
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 11790 20040 11796 20052
rect 11379 20012 11796 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 12618 20000 12624 20052
rect 12676 20000 12682 20052
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 13909 20043 13967 20049
rect 13909 20040 13921 20043
rect 13872 20012 13921 20040
rect 13872 20000 13878 20012
rect 13909 20009 13921 20012
rect 13955 20009 13967 20043
rect 13909 20003 13967 20009
rect 12526 19972 12532 19984
rect 10181 19876 10548 19904
rect 11072 19944 12532 19972
rect 10181 19873 10193 19876
rect 10135 19867 10193 19873
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19805 7435 19839
rect 7711 19839 7769 19845
rect 7711 19836 7723 19839
rect 7377 19799 7435 19805
rect 7484 19808 7723 19836
rect 6087 19789 6145 19795
rect 6104 19700 6132 19789
rect 6932 19768 6960 19796
rect 7484 19768 7512 19808
rect 7711 19805 7723 19808
rect 7757 19836 7769 19839
rect 8202 19836 8208 19848
rect 7757 19808 8208 19836
rect 7757 19805 7769 19808
rect 7711 19799 7769 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 9950 19796 9956 19848
rect 10008 19845 10014 19848
rect 11072 19845 11100 19944
rect 12526 19932 12532 19944
rect 12584 19932 12590 19984
rect 12636 19972 12664 20000
rect 12713 19975 12771 19981
rect 12713 19972 12725 19975
rect 12636 19944 12725 19972
rect 12713 19941 12725 19944
rect 12759 19941 12771 19975
rect 12713 19935 12771 19941
rect 11330 19864 11336 19916
rect 11388 19904 11394 19916
rect 12069 19907 12127 19913
rect 12069 19904 12081 19907
rect 11388 19876 12081 19904
rect 11388 19864 11394 19876
rect 12069 19873 12081 19876
rect 12115 19904 12127 19907
rect 12342 19904 12348 19916
rect 12115 19876 12348 19904
rect 12115 19873 12127 19876
rect 12069 19867 12127 19873
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 12989 19907 13047 19913
rect 12989 19904 13001 19907
rect 12860 19876 13001 19904
rect 12860 19864 12866 19876
rect 12989 19873 13001 19876
rect 13035 19873 13047 19907
rect 12989 19867 13047 19873
rect 13127 19907 13185 19913
rect 13127 19873 13139 19907
rect 13173 19904 13185 19907
rect 13446 19904 13452 19916
rect 13173 19876 13452 19904
rect 13173 19873 13185 19876
rect 13127 19867 13185 19873
rect 13446 19864 13452 19876
rect 13504 19904 13510 19916
rect 13630 19904 13636 19916
rect 13504 19876 13636 19904
rect 13504 19864 13510 19876
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 10008 19839 10036 19845
rect 10024 19805 10036 19839
rect 10008 19799 10036 19805
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19805 11115 19839
rect 12253 19839 12311 19845
rect 12253 19836 12265 19839
rect 11057 19799 11115 19805
rect 11164 19808 12265 19836
rect 10008 19796 10014 19799
rect 6932 19740 7512 19768
rect 10686 19728 10692 19780
rect 10744 19768 10750 19780
rect 11164 19768 11192 19808
rect 12253 19805 12265 19808
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 13262 19796 13268 19848
rect 13320 19796 13326 19848
rect 10744 19740 11192 19768
rect 11609 19771 11667 19777
rect 10744 19728 10750 19740
rect 11609 19737 11621 19771
rect 11655 19737 11667 19771
rect 11609 19731 11667 19737
rect 11977 19771 12035 19777
rect 11977 19737 11989 19771
rect 12023 19737 12035 19771
rect 11977 19731 12035 19737
rect 1176 19672 6132 19700
rect 1176 19660 1182 19672
rect 7190 19660 7196 19712
rect 7248 19660 7254 19712
rect 9306 19660 9312 19712
rect 9364 19700 9370 19712
rect 11624 19700 11652 19731
rect 9364 19672 11652 19700
rect 11992 19700 12020 19731
rect 15194 19728 15200 19780
rect 15252 19768 15258 19780
rect 15470 19768 15476 19780
rect 15252 19740 15476 19768
rect 15252 19728 15258 19740
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 13814 19700 13820 19712
rect 11992 19672 13820 19700
rect 9364 19660 9370 19672
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 1104 19610 14971 19632
rect 1104 19558 4376 19610
rect 4428 19558 4440 19610
rect 4492 19558 4504 19610
rect 4556 19558 4568 19610
rect 4620 19558 4632 19610
rect 4684 19558 7803 19610
rect 7855 19558 7867 19610
rect 7919 19558 7931 19610
rect 7983 19558 7995 19610
rect 8047 19558 8059 19610
rect 8111 19558 11230 19610
rect 11282 19558 11294 19610
rect 11346 19558 11358 19610
rect 11410 19558 11422 19610
rect 11474 19558 11486 19610
rect 11538 19558 14657 19610
rect 14709 19558 14721 19610
rect 14773 19558 14785 19610
rect 14837 19558 14849 19610
rect 14901 19558 14913 19610
rect 14965 19558 14971 19610
rect 1104 19536 14971 19558
rect 7098 19456 7104 19508
rect 7156 19456 7162 19508
rect 7190 19456 7196 19508
rect 7248 19456 7254 19508
rect 7392 19468 7696 19496
rect 6730 19388 6736 19440
rect 6788 19428 6794 19440
rect 6788 19400 7052 19428
rect 6788 19388 6794 19400
rect 1486 19320 1492 19372
rect 1544 19320 1550 19372
rect 6822 19320 6828 19372
rect 6880 19320 6886 19372
rect 7024 19369 7052 19400
rect 7116 19369 7144 19456
rect 7208 19428 7236 19456
rect 7392 19437 7420 19468
rect 7377 19431 7435 19437
rect 7208 19400 7328 19428
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19329 7067 19363
rect 7009 19323 7067 19329
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19329 7159 19363
rect 7300 19360 7328 19400
rect 7377 19397 7389 19431
rect 7423 19397 7435 19431
rect 7668 19428 7696 19468
rect 7742 19456 7748 19508
rect 7800 19496 7806 19508
rect 9030 19496 9036 19508
rect 7800 19468 9036 19496
rect 7800 19456 7806 19468
rect 9030 19456 9036 19468
rect 9088 19496 9094 19508
rect 9088 19468 10824 19496
rect 9088 19456 9094 19468
rect 10796 19428 10824 19468
rect 10870 19456 10876 19508
rect 10928 19496 10934 19508
rect 11057 19499 11115 19505
rect 11057 19496 11069 19499
rect 10928 19468 11069 19496
rect 10928 19456 10934 19468
rect 11057 19465 11069 19468
rect 11103 19465 11115 19499
rect 11057 19459 11115 19465
rect 11146 19456 11152 19508
rect 11204 19456 11210 19508
rect 12526 19456 12532 19508
rect 12584 19496 12590 19508
rect 12584 19468 13216 19496
rect 12584 19456 12590 19468
rect 11164 19428 11192 19456
rect 7668 19400 10732 19428
rect 10796 19400 11008 19428
rect 11164 19400 11560 19428
rect 7377 19391 7435 19397
rect 7469 19363 7527 19369
rect 7469 19360 7481 19363
rect 7300 19332 7481 19360
rect 7101 19323 7159 19329
rect 7469 19329 7481 19332
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 7558 19320 7564 19372
rect 7616 19320 7622 19372
rect 8202 19360 8208 19372
rect 8163 19332 8208 19360
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 10318 19320 10324 19372
rect 10376 19360 10382 19372
rect 10594 19360 10600 19372
rect 10376 19332 10600 19360
rect 10376 19320 10382 19332
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 6917 19295 6975 19301
rect 6917 19261 6929 19295
rect 6963 19292 6975 19295
rect 7190 19292 7196 19315
rect 6963 19264 7196 19292
rect 6963 19261 6975 19264
rect 7190 19263 7196 19264
rect 7248 19263 7254 19315
rect 6917 19255 6975 19261
rect 7374 19252 7380 19304
rect 7432 19292 7438 19304
rect 7576 19292 7604 19320
rect 7929 19295 7987 19301
rect 7929 19292 7941 19295
rect 7432 19264 7477 19292
rect 7576 19264 7941 19292
rect 7432 19252 7438 19264
rect 7929 19261 7941 19264
rect 7975 19261 7987 19295
rect 10704 19292 10732 19400
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19360 10839 19363
rect 10870 19360 10876 19372
rect 10827 19332 10876 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 10980 19360 11008 19400
rect 11532 19369 11560 19400
rect 11241 19363 11299 19369
rect 11241 19360 11253 19363
rect 10980 19332 11253 19360
rect 11241 19329 11253 19332
rect 11287 19329 11299 19363
rect 11241 19323 11299 19329
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19329 11575 19363
rect 12069 19363 12127 19369
rect 12069 19360 12081 19363
rect 11517 19323 11575 19329
rect 11624 19332 12081 19360
rect 11624 19292 11652 19332
rect 12069 19329 12081 19332
rect 12115 19329 12127 19363
rect 12069 19323 12127 19329
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 12713 19363 12771 19369
rect 12713 19360 12725 19363
rect 12308 19332 12725 19360
rect 12308 19320 12314 19332
rect 10704 19264 11652 19292
rect 7929 19255 7987 19261
rect 1673 19227 1731 19233
rect 1673 19193 1685 19227
rect 1719 19224 1731 19227
rect 3510 19224 3516 19236
rect 1719 19196 3516 19224
rect 1719 19193 1731 19196
rect 1673 19187 1731 19193
rect 3510 19184 3516 19196
rect 3568 19184 3574 19236
rect 7193 19227 7251 19233
rect 3620 19196 7144 19224
rect 3620 19168 3648 19196
rect 3602 19116 3608 19168
rect 3660 19116 3666 19168
rect 5718 19116 5724 19168
rect 5776 19156 5782 19168
rect 5994 19156 6000 19168
rect 5776 19128 6000 19156
rect 5776 19116 5782 19128
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 7116 19156 7144 19196
rect 7193 19193 7205 19227
rect 7239 19224 7251 19227
rect 7561 19227 7619 19233
rect 7561 19224 7573 19227
rect 7239 19196 7573 19224
rect 7239 19193 7251 19196
rect 7193 19187 7251 19193
rect 7561 19193 7573 19196
rect 7607 19193 7619 19227
rect 7561 19187 7619 19193
rect 7650 19156 7656 19168
rect 7116 19128 7656 19156
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 7944 19156 7972 19255
rect 11698 19252 11704 19304
rect 11756 19292 11762 19304
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 11756 19264 11805 19292
rect 11756 19252 11762 19264
rect 11793 19261 11805 19264
rect 11839 19261 11851 19295
rect 12544 19292 12572 19332
rect 12713 19329 12725 19332
rect 12759 19329 12771 19363
rect 12713 19323 12771 19329
rect 12955 19363 13013 19369
rect 12955 19329 12967 19363
rect 13001 19360 13013 19363
rect 13078 19360 13084 19372
rect 13001 19332 13084 19360
rect 13001 19329 13013 19332
rect 12955 19323 13013 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 13188 19360 13216 19468
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13725 19499 13783 19505
rect 13725 19496 13737 19499
rect 13320 19468 13737 19496
rect 13320 19456 13326 19468
rect 13725 19465 13737 19468
rect 13771 19465 13783 19499
rect 13725 19459 13783 19465
rect 14366 19456 14372 19508
rect 14424 19456 14430 19508
rect 14458 19456 14464 19508
rect 14516 19496 14522 19508
rect 14642 19496 14648 19508
rect 14516 19468 14648 19496
rect 14516 19456 14522 19468
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 14185 19363 14243 19369
rect 13188 19332 13860 19360
rect 13832 19304 13860 19332
rect 14185 19329 14197 19363
rect 14231 19360 14243 19363
rect 14458 19360 14464 19372
rect 14231 19332 14464 19360
rect 14231 19329 14243 19332
rect 14185 19323 14243 19329
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 11793 19255 11851 19261
rect 12268 19264 12572 19292
rect 9398 19224 9404 19236
rect 8864 19196 9404 19224
rect 8864 19156 8892 19196
rect 9398 19184 9404 19196
rect 9456 19184 9462 19236
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10686 19224 10692 19236
rect 10008 19196 10692 19224
rect 10008 19184 10014 19196
rect 10686 19184 10692 19196
rect 10744 19184 10750 19236
rect 10873 19227 10931 19233
rect 10873 19193 10885 19227
rect 10919 19224 10931 19227
rect 11609 19227 11667 19233
rect 11609 19224 11621 19227
rect 10919 19196 11621 19224
rect 10919 19193 10931 19196
rect 10873 19187 10931 19193
rect 11609 19193 11621 19196
rect 11655 19193 11667 19227
rect 11609 19187 11667 19193
rect 12268 19168 12296 19264
rect 13814 19252 13820 19304
rect 13872 19252 13878 19304
rect 7944 19128 8892 19156
rect 8938 19116 8944 19168
rect 8996 19116 9002 19168
rect 11698 19116 11704 19168
rect 11756 19116 11762 19168
rect 12250 19116 12256 19168
rect 12308 19116 12314 19168
rect 12345 19159 12403 19165
rect 12345 19125 12357 19159
rect 12391 19156 12403 19159
rect 14090 19156 14096 19168
rect 12391 19128 14096 19156
rect 12391 19125 12403 19128
rect 12345 19119 12403 19125
rect 14090 19116 14096 19128
rect 14148 19116 14154 19168
rect 1104 19066 14812 19088
rect 1104 19014 2663 19066
rect 2715 19014 2727 19066
rect 2779 19014 2791 19066
rect 2843 19014 2855 19066
rect 2907 19014 2919 19066
rect 2971 19014 6090 19066
rect 6142 19014 6154 19066
rect 6206 19014 6218 19066
rect 6270 19014 6282 19066
rect 6334 19014 6346 19066
rect 6398 19014 9517 19066
rect 9569 19014 9581 19066
rect 9633 19014 9645 19066
rect 9697 19014 9709 19066
rect 9761 19014 9773 19066
rect 9825 19014 12944 19066
rect 12996 19014 13008 19066
rect 13060 19014 13072 19066
rect 13124 19014 13136 19066
rect 13188 19014 13200 19066
rect 13252 19014 14812 19066
rect 1104 18992 14812 19014
rect 3878 18912 3884 18964
rect 3936 18952 3942 18964
rect 4706 18952 4712 18964
rect 3936 18924 4712 18952
rect 3936 18912 3942 18924
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 5261 18955 5319 18961
rect 5261 18921 5273 18955
rect 5307 18952 5319 18955
rect 8754 18952 8760 18964
rect 5307 18924 8760 18952
rect 5307 18921 5319 18924
rect 5261 18915 5319 18921
rect 8754 18912 8760 18924
rect 8812 18952 8818 18964
rect 11885 18955 11943 18961
rect 8812 18924 10548 18952
rect 8812 18912 8818 18924
rect 6457 18887 6515 18893
rect 6457 18853 6469 18887
rect 6503 18884 6515 18887
rect 6914 18884 6920 18896
rect 6503 18856 6920 18884
rect 6503 18853 6515 18856
rect 6457 18847 6515 18853
rect 6914 18844 6920 18856
rect 6972 18844 6978 18896
rect 7190 18884 7196 18896
rect 7116 18856 7196 18884
rect 6932 18816 6960 18844
rect 7116 18825 7144 18856
rect 7190 18844 7196 18856
rect 7248 18844 7254 18896
rect 7285 18887 7343 18893
rect 7285 18853 7297 18887
rect 7331 18853 7343 18887
rect 7285 18847 7343 18853
rect 6840 18788 6960 18816
rect 7101 18819 7159 18825
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18717 5503 18751
rect 5445 18711 5503 18717
rect 3970 18640 3976 18692
rect 4028 18680 4034 18692
rect 5169 18683 5227 18689
rect 5169 18680 5181 18683
rect 4028 18652 5181 18680
rect 4028 18640 4034 18652
rect 5169 18649 5181 18652
rect 5215 18649 5227 18683
rect 5460 18680 5488 18711
rect 5626 18708 5632 18760
rect 5684 18748 5690 18760
rect 6840 18757 6868 18788
rect 7101 18785 7113 18819
rect 7147 18785 7159 18819
rect 7300 18816 7328 18847
rect 7650 18844 7656 18896
rect 7708 18844 7714 18896
rect 7834 18844 7840 18896
rect 7892 18884 7898 18896
rect 9674 18884 9680 18896
rect 7892 18856 9680 18884
rect 7892 18844 7898 18856
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 7300 18788 7604 18816
rect 7101 18779 7159 18785
rect 5719 18751 5777 18757
rect 5719 18748 5731 18751
rect 5684 18720 5731 18748
rect 5684 18708 5690 18720
rect 5719 18717 5731 18720
rect 5765 18748 5777 18751
rect 6825 18751 6883 18757
rect 5765 18720 6776 18748
rect 5765 18717 5777 18720
rect 5719 18711 5777 18717
rect 5810 18680 5816 18692
rect 5460 18652 5816 18680
rect 5169 18643 5227 18649
rect 5810 18640 5816 18652
rect 5868 18680 5874 18692
rect 5994 18680 6000 18692
rect 5868 18652 6000 18680
rect 5868 18640 5874 18652
rect 5994 18640 6000 18652
rect 6052 18640 6058 18692
rect 6748 18624 6776 18720
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 6917 18751 6975 18757
rect 6917 18717 6929 18751
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 6932 18680 6960 18711
rect 7374 18708 7380 18760
rect 7432 18748 7438 18760
rect 7576 18757 7604 18788
rect 7469 18751 7527 18757
rect 7469 18748 7481 18751
rect 7432 18720 7481 18748
rect 7432 18708 7438 18720
rect 7469 18717 7481 18720
rect 7515 18717 7527 18751
rect 7469 18711 7527 18717
rect 7561 18751 7619 18757
rect 7561 18717 7573 18751
rect 7607 18717 7619 18751
rect 7668 18748 7696 18844
rect 7668 18720 8524 18748
rect 7561 18711 7619 18717
rect 7653 18683 7711 18689
rect 7653 18680 7665 18683
rect 6932 18652 7665 18680
rect 7653 18649 7665 18652
rect 7699 18649 7711 18683
rect 8496 18680 8524 18720
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 9858 18748 9864 18760
rect 8628 18720 9864 18748
rect 8628 18708 8634 18720
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 10520 18748 10548 18924
rect 11885 18921 11897 18955
rect 11931 18952 11943 18955
rect 11974 18952 11980 18964
rect 11931 18924 11980 18952
rect 11931 18921 11943 18924
rect 11885 18915 11943 18921
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 12437 18955 12495 18961
rect 12437 18921 12449 18955
rect 12483 18952 12495 18955
rect 14274 18952 14280 18964
rect 12483 18924 14280 18952
rect 12483 18921 12495 18924
rect 12437 18915 12495 18921
rect 14274 18912 14280 18924
rect 14332 18912 14338 18964
rect 11606 18776 11612 18828
rect 11664 18776 11670 18828
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 11756 18788 12204 18816
rect 11756 18776 11762 18788
rect 11425 18751 11483 18757
rect 11425 18748 11437 18751
rect 10119 18721 10177 18727
rect 10119 18718 10131 18721
rect 10060 18690 10131 18718
rect 10060 18680 10088 18690
rect 10119 18687 10131 18690
rect 10165 18687 10177 18721
rect 10520 18720 11437 18748
rect 11425 18717 11437 18720
rect 11471 18717 11483 18751
rect 11624 18748 11652 18776
rect 12176 18757 12204 18788
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 12621 18819 12679 18825
rect 12621 18816 12633 18819
rect 12308 18788 12633 18816
rect 12308 18776 12314 18788
rect 12360 18760 12388 18788
rect 12621 18785 12633 18788
rect 12667 18785 12679 18819
rect 12621 18779 12679 18785
rect 11425 18711 11483 18717
rect 11532 18720 11652 18748
rect 12161 18751 12219 18757
rect 10119 18681 10177 18687
rect 8496 18652 10088 18680
rect 7653 18643 7711 18649
rect 10318 18640 10324 18692
rect 10376 18680 10382 18692
rect 11532 18680 11560 18720
rect 12161 18717 12173 18751
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 12342 18708 12348 18760
rect 12400 18708 12406 18760
rect 12863 18751 12921 18757
rect 12863 18717 12875 18751
rect 12909 18748 12921 18751
rect 12986 18748 12992 18760
rect 12909 18720 12992 18748
rect 12909 18717 12921 18720
rect 12863 18711 12921 18717
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 13998 18748 14004 18760
rect 13872 18720 14004 18748
rect 13872 18708 13878 18720
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 14550 18748 14556 18760
rect 14323 18720 14556 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 10376 18652 11560 18680
rect 10376 18640 10382 18652
rect 11606 18640 11612 18692
rect 11664 18640 11670 18692
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 14292 18680 14320 18711
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 12308 18652 14320 18680
rect 12308 18640 12314 18652
rect 6730 18572 6736 18624
rect 6788 18572 6794 18624
rect 7098 18572 7104 18624
rect 7156 18572 7162 18624
rect 10870 18572 10876 18624
rect 10928 18572 10934 18624
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 11241 18615 11299 18621
rect 11241 18612 11253 18615
rect 11204 18584 11253 18612
rect 11204 18572 11210 18584
rect 11241 18581 11253 18584
rect 11287 18581 11299 18615
rect 11241 18575 11299 18581
rect 11882 18572 11888 18624
rect 11940 18612 11946 18624
rect 13538 18612 13544 18624
rect 11940 18584 13544 18612
rect 11940 18572 11946 18584
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 13633 18615 13691 18621
rect 13633 18581 13645 18615
rect 13679 18612 13691 18615
rect 13814 18612 13820 18624
rect 13679 18584 13820 18612
rect 13679 18581 13691 18584
rect 13633 18575 13691 18581
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 14090 18572 14096 18624
rect 14148 18572 14154 18624
rect 1104 18522 14971 18544
rect 1104 18470 4376 18522
rect 4428 18470 4440 18522
rect 4492 18470 4504 18522
rect 4556 18470 4568 18522
rect 4620 18470 4632 18522
rect 4684 18470 7803 18522
rect 7855 18470 7867 18522
rect 7919 18470 7931 18522
rect 7983 18470 7995 18522
rect 8047 18470 8059 18522
rect 8111 18470 11230 18522
rect 11282 18470 11294 18522
rect 11346 18470 11358 18522
rect 11410 18470 11422 18522
rect 11474 18470 11486 18522
rect 11538 18470 14657 18522
rect 14709 18470 14721 18522
rect 14773 18470 14785 18522
rect 14837 18470 14849 18522
rect 14901 18470 14913 18522
rect 14965 18470 14971 18522
rect 1104 18448 14971 18470
rect 6822 18368 6828 18420
rect 6880 18368 6886 18420
rect 10870 18368 10876 18420
rect 10928 18368 10934 18420
rect 11146 18368 11152 18420
rect 11204 18368 11210 18420
rect 11333 18411 11391 18417
rect 11333 18377 11345 18411
rect 11379 18408 11391 18411
rect 11882 18408 11888 18420
rect 11379 18380 11888 18408
rect 11379 18377 11391 18380
rect 11333 18371 11391 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 14090 18408 14096 18420
rect 12268 18380 14096 18408
rect 8662 18340 8668 18352
rect 2746 18312 8668 18340
rect 750 18232 756 18284
rect 808 18272 814 18284
rect 1489 18275 1547 18281
rect 1489 18272 1501 18275
rect 808 18244 1501 18272
rect 808 18232 814 18244
rect 1489 18241 1501 18244
rect 1535 18241 1547 18275
rect 1489 18235 1547 18241
rect 1673 18139 1731 18145
rect 1673 18105 1685 18139
rect 1719 18105 1731 18139
rect 1673 18099 1731 18105
rect 1688 18068 1716 18099
rect 2746 18068 2774 18312
rect 8662 18300 8668 18312
rect 8720 18300 8726 18352
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 5057 18275 5115 18281
rect 5057 18272 5069 18275
rect 4028 18244 5069 18272
rect 4028 18232 4034 18244
rect 5057 18241 5069 18244
rect 5103 18241 5115 18275
rect 5057 18235 5115 18241
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18272 7067 18275
rect 7466 18272 7472 18284
rect 7055 18244 7472 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 4246 18164 4252 18216
rect 4304 18204 4310 18216
rect 4798 18204 4804 18216
rect 4304 18176 4804 18204
rect 4304 18164 4310 18176
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 5810 18164 5816 18216
rect 5868 18204 5874 18216
rect 6638 18204 6644 18216
rect 5868 18176 6644 18204
rect 5868 18164 5874 18176
rect 6638 18164 6644 18176
rect 6696 18164 6702 18216
rect 6181 18139 6239 18145
rect 6181 18105 6193 18139
rect 6227 18136 6239 18139
rect 7024 18136 7052 18235
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 8815 18275 8873 18281
rect 8815 18272 8827 18275
rect 8496 18244 8827 18272
rect 6227 18108 7052 18136
rect 6227 18105 6239 18108
rect 6181 18099 6239 18105
rect 7466 18096 7472 18148
rect 7524 18136 7530 18148
rect 8496 18136 8524 18244
rect 8815 18241 8827 18244
rect 8861 18272 8873 18275
rect 9582 18272 9588 18284
rect 8861 18244 9588 18272
rect 8861 18241 8873 18244
rect 8815 18235 8873 18241
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18173 8631 18207
rect 8573 18167 8631 18173
rect 7524 18108 8524 18136
rect 7524 18096 7530 18108
rect 8588 18080 8616 18167
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 10134 18204 10140 18216
rect 9456 18176 10140 18204
rect 9456 18164 9462 18176
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 10888 18204 10916 18368
rect 11164 18340 11192 18368
rect 11164 18312 12204 18340
rect 11146 18232 11152 18284
rect 11204 18232 11210 18284
rect 12176 18281 12204 18312
rect 12268 18281 12296 18380
rect 14090 18368 14096 18380
rect 14148 18368 14154 18420
rect 14458 18368 14464 18420
rect 14516 18368 14522 18420
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 11977 18275 12035 18281
rect 11977 18272 11989 18275
rect 11563 18244 11989 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11977 18241 11989 18244
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 12161 18275 12219 18281
rect 12161 18241 12173 18275
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 11532 18204 11560 18235
rect 13814 18232 13820 18284
rect 13872 18232 13878 18284
rect 10888 18176 11560 18204
rect 11793 18207 11851 18213
rect 11793 18173 11805 18207
rect 11839 18204 11851 18207
rect 12069 18207 12127 18213
rect 12069 18204 12081 18207
rect 11839 18176 12081 18204
rect 11839 18173 11851 18176
rect 11793 18167 11851 18173
rect 12069 18173 12081 18176
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 12526 18164 12532 18216
rect 12584 18204 12590 18216
rect 12621 18207 12679 18213
rect 12621 18204 12633 18207
rect 12584 18176 12633 18204
rect 12584 18164 12590 18176
rect 12621 18173 12633 18176
rect 12667 18173 12679 18207
rect 12621 18167 12679 18173
rect 12710 18164 12716 18216
rect 12768 18164 12774 18216
rect 12802 18164 12808 18216
rect 12860 18164 12866 18216
rect 13541 18207 13599 18213
rect 13541 18204 13553 18207
rect 13121 18176 13553 18204
rect 11609 18139 11667 18145
rect 11609 18105 11621 18139
rect 11655 18136 11667 18139
rect 12345 18139 12403 18145
rect 12345 18136 12357 18139
rect 11655 18108 12357 18136
rect 11655 18105 11667 18108
rect 11609 18099 11667 18105
rect 12345 18105 12357 18108
rect 12391 18105 12403 18139
rect 12728 18136 12756 18164
rect 13121 18136 13149 18176
rect 13541 18173 13553 18176
rect 13587 18173 13599 18207
rect 13541 18167 13599 18173
rect 13630 18164 13636 18216
rect 13688 18213 13694 18216
rect 13688 18207 13716 18213
rect 13704 18173 13716 18207
rect 13688 18167 13716 18173
rect 13688 18164 13694 18167
rect 12728 18108 13149 18136
rect 12345 18099 12403 18105
rect 13262 18096 13268 18148
rect 13320 18096 13326 18148
rect 1688 18040 2774 18068
rect 5994 18028 6000 18080
rect 6052 18068 6058 18080
rect 8570 18068 8576 18080
rect 6052 18040 8576 18068
rect 6052 18028 6058 18040
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 9398 18028 9404 18080
rect 9456 18068 9462 18080
rect 9585 18071 9643 18077
rect 9585 18068 9597 18071
rect 9456 18040 9597 18068
rect 9456 18028 9462 18040
rect 9585 18037 9597 18040
rect 9631 18037 9643 18071
rect 9585 18031 9643 18037
rect 11701 18071 11759 18077
rect 11701 18037 11713 18071
rect 11747 18068 11759 18071
rect 13354 18068 13360 18080
rect 11747 18040 13360 18068
rect 11747 18037 11759 18040
rect 11701 18031 11759 18037
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14458 18068 14464 18080
rect 13872 18040 14464 18068
rect 13872 18028 13878 18040
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 1104 17978 14812 18000
rect 1104 17926 2663 17978
rect 2715 17926 2727 17978
rect 2779 17926 2791 17978
rect 2843 17926 2855 17978
rect 2907 17926 2919 17978
rect 2971 17926 6090 17978
rect 6142 17926 6154 17978
rect 6206 17926 6218 17978
rect 6270 17926 6282 17978
rect 6334 17926 6346 17978
rect 6398 17926 9517 17978
rect 9569 17926 9581 17978
rect 9633 17926 9645 17978
rect 9697 17926 9709 17978
rect 9761 17926 9773 17978
rect 9825 17926 12944 17978
rect 12996 17926 13008 17978
rect 13060 17926 13072 17978
rect 13124 17926 13136 17978
rect 13188 17926 13200 17978
rect 13252 17926 14812 17978
rect 1104 17904 14812 17926
rect 7006 17824 7012 17876
rect 7064 17864 7070 17876
rect 7558 17864 7564 17876
rect 7064 17836 7564 17864
rect 7064 17824 7070 17836
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 9214 17864 9220 17876
rect 8444 17836 9220 17864
rect 8444 17824 8450 17836
rect 9214 17824 9220 17836
rect 9272 17864 9278 17876
rect 9272 17836 10640 17864
rect 9272 17824 9278 17836
rect 1673 17799 1731 17805
rect 1673 17765 1685 17799
rect 1719 17796 1731 17799
rect 5810 17796 5816 17808
rect 1719 17768 5816 17796
rect 1719 17765 1731 17768
rect 1673 17759 1731 17765
rect 5810 17756 5816 17768
rect 5868 17756 5874 17808
rect 10612 17796 10640 17836
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 11609 17867 11667 17873
rect 11609 17864 11621 17867
rect 10744 17836 11621 17864
rect 10744 17824 10750 17836
rect 11609 17833 11621 17836
rect 11655 17833 11667 17867
rect 11609 17827 11667 17833
rect 11698 17824 11704 17876
rect 11756 17864 11762 17876
rect 11885 17867 11943 17873
rect 11885 17864 11897 17867
rect 11756 17836 11897 17864
rect 11756 17824 11762 17836
rect 11885 17833 11897 17836
rect 11931 17833 11943 17867
rect 11885 17827 11943 17833
rect 13262 17824 13268 17876
rect 13320 17824 13326 17876
rect 13814 17824 13820 17876
rect 13872 17824 13878 17876
rect 10870 17796 10876 17808
rect 10612 17768 10876 17796
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 11333 17799 11391 17805
rect 11333 17765 11345 17799
rect 11379 17796 11391 17799
rect 11379 17768 12112 17796
rect 11379 17765 11391 17768
rect 11333 17759 11391 17765
rect 12084 17740 12112 17768
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 8628 17700 9413 17728
rect 8628 17688 8634 17700
rect 9401 17697 9413 17700
rect 9447 17697 9459 17731
rect 11698 17728 11704 17740
rect 9401 17691 9459 17697
rect 11164 17700 11704 17728
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 6181 17663 6239 17669
rect 6181 17660 6193 17663
rect 6052 17632 6193 17660
rect 6052 17620 6058 17632
rect 6181 17629 6193 17632
rect 6227 17629 6239 17663
rect 6181 17623 6239 17629
rect 6439 17633 6497 17639
rect 750 17552 756 17604
rect 808 17592 814 17604
rect 1489 17595 1547 17601
rect 1489 17592 1501 17595
rect 808 17564 1501 17592
rect 808 17552 814 17564
rect 1489 17561 1501 17564
rect 1535 17561 1547 17595
rect 6439 17599 6451 17633
rect 6485 17630 6497 17633
rect 6485 17604 6500 17630
rect 7098 17620 7104 17672
rect 7156 17620 7162 17672
rect 9674 17660 9680 17672
rect 9635 17632 9680 17660
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 11164 17669 11192 17700
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 12066 17688 12072 17740
rect 12124 17688 12130 17740
rect 13538 17688 13544 17740
rect 13596 17728 13602 17740
rect 14642 17728 14648 17740
rect 13596 17700 14648 17728
rect 13596 17688 13602 17700
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 11422 17620 11428 17672
rect 11480 17620 11486 17672
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 12253 17663 12311 17669
rect 12253 17660 12265 17663
rect 11572 17632 12265 17660
rect 11572 17620 11578 17632
rect 12253 17629 12265 17632
rect 12299 17629 12311 17663
rect 12253 17623 12311 17629
rect 12495 17663 12553 17669
rect 12495 17629 12507 17663
rect 12541 17660 12553 17663
rect 13633 17663 13691 17669
rect 12541 17629 12554 17660
rect 12495 17623 12554 17629
rect 13633 17629 13645 17663
rect 13679 17660 13691 17663
rect 15194 17660 15200 17672
rect 13679 17632 15200 17660
rect 13679 17629 13691 17632
rect 13633 17623 13691 17629
rect 6439 17593 6460 17599
rect 1489 17555 1547 17561
rect 6454 17552 6460 17593
rect 6512 17552 6518 17604
rect 7116 17592 7144 17620
rect 11793 17595 11851 17601
rect 11793 17592 11805 17595
rect 7116 17564 11805 17592
rect 11793 17561 11805 17564
rect 11839 17561 11851 17595
rect 12268 17592 12296 17623
rect 12342 17592 12348 17604
rect 12268 17564 12348 17592
rect 11793 17555 11851 17561
rect 12342 17552 12348 17564
rect 12400 17552 12406 17604
rect 3602 17484 3608 17536
rect 3660 17524 3666 17536
rect 6472 17524 6500 17552
rect 3660 17496 6500 17524
rect 3660 17484 3666 17496
rect 7190 17484 7196 17536
rect 7248 17484 7254 17536
rect 10413 17527 10471 17533
rect 10413 17493 10425 17527
rect 10459 17524 10471 17527
rect 10686 17524 10692 17536
rect 10459 17496 10692 17524
rect 10459 17493 10471 17496
rect 10413 17487 10471 17493
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 12526 17524 12554 17623
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 10928 17496 12554 17524
rect 10928 17484 10934 17496
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 15194 17348 15200 17400
rect 15252 17388 15258 17400
rect 15930 17388 15936 17400
rect 15252 17360 15936 17388
rect 15252 17348 15258 17360
rect 15930 17348 15936 17360
rect 15988 17348 15994 17400
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 1670 17320 1676 17332
rect 1627 17292 1676 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 7190 17280 7196 17332
rect 7248 17280 7254 17332
rect 8941 17323 8999 17329
rect 8941 17289 8953 17323
rect 8987 17320 8999 17323
rect 9306 17320 9312 17332
rect 8987 17292 9312 17320
rect 8987 17289 8999 17292
rect 8941 17283 8999 17289
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 11379 17292 11834 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 1486 17144 1492 17196
rect 1544 17144 1550 17196
rect 7006 17144 7012 17196
rect 7064 17184 7070 17196
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 7064 17156 7113 17184
rect 7064 17144 7070 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 7208 17184 7236 17280
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11806 17252 11834 17292
rect 12618 17280 12624 17332
rect 12676 17320 12682 17332
rect 13265 17323 13323 17329
rect 13265 17320 13277 17323
rect 12676 17292 13277 17320
rect 12676 17280 12682 17292
rect 13265 17289 13277 17292
rect 13311 17320 13323 17323
rect 13630 17320 13636 17332
rect 13311 17292 13636 17320
rect 13311 17289 13323 17292
rect 13265 17283 13323 17289
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 13817 17323 13875 17329
rect 13817 17289 13829 17323
rect 13863 17320 13875 17323
rect 13906 17320 13912 17332
rect 13863 17292 13912 17320
rect 13863 17289 13875 17292
rect 13817 17283 13875 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14369 17323 14427 17329
rect 14369 17289 14381 17323
rect 14415 17320 14427 17323
rect 15470 17320 15476 17332
rect 14415 17292 15476 17320
rect 14415 17289 14427 17292
rect 14369 17283 14427 17289
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 14093 17255 14151 17261
rect 14093 17252 14105 17255
rect 11480 17224 11742 17252
rect 11806 17224 14105 17252
rect 11480 17212 11486 17224
rect 8202 17193 8208 17196
rect 8159 17187 8208 17193
rect 7208 17156 7512 17184
rect 7101 17147 7159 17153
rect 1394 17076 1400 17128
rect 1452 17116 1458 17128
rect 1670 17116 1676 17128
rect 1452 17088 1676 17116
rect 1452 17076 1458 17088
rect 1670 17076 1676 17088
rect 1728 17076 1734 17128
rect 7282 17076 7288 17128
rect 7340 17076 7346 17128
rect 7484 17116 7512 17156
rect 8159 17153 8171 17187
rect 8205 17153 8208 17187
rect 8159 17147 8208 17153
rect 8202 17144 8208 17147
rect 8260 17144 8266 17196
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 9858 17184 9864 17196
rect 9539 17156 9864 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 10410 17144 10416 17196
rect 10468 17144 10474 17196
rect 10686 17144 10692 17196
rect 10744 17144 10750 17196
rect 11714 17184 11742 17224
rect 14093 17221 14105 17224
rect 14139 17221 14151 17255
rect 14093 17215 14151 17221
rect 11851 17187 11909 17193
rect 11851 17184 11863 17187
rect 11714 17156 11863 17184
rect 11851 17153 11863 17156
rect 11897 17153 11909 17187
rect 11851 17147 11909 17153
rect 13170 17144 13176 17196
rect 13228 17144 13234 17196
rect 13354 17144 13360 17196
rect 13412 17184 13418 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 13412 17156 13553 17184
rect 13412 17144 13418 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7484 17088 7757 17116
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7745 17079 7803 17085
rect 7852 17088 8033 17116
rect 7852 16980 7880 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 8294 17076 8300 17128
rect 8352 17076 8358 17128
rect 9398 17076 9404 17128
rect 9456 17076 9462 17128
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17116 9735 17119
rect 10551 17119 10609 17125
rect 9723 17088 10272 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 9416 17048 9444 17076
rect 10137 17051 10195 17057
rect 10137 17048 10149 17051
rect 9416 17020 10149 17048
rect 10137 17017 10149 17020
rect 10183 17017 10195 17051
rect 10137 17011 10195 17017
rect 10042 16980 10048 16992
rect 7852 16952 10048 16980
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10244 16980 10272 17088
rect 10551 17085 10563 17119
rect 10597 17116 10609 17119
rect 10870 17116 10876 17128
rect 10597 17088 10876 17116
rect 10597 17085 10609 17088
rect 10551 17079 10609 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 11238 17076 11244 17128
rect 11296 17116 11302 17128
rect 11609 17119 11667 17125
rect 11609 17116 11621 17119
rect 11296 17088 11621 17116
rect 11296 17076 11302 17088
rect 11609 17085 11621 17088
rect 11655 17085 11667 17119
rect 11609 17079 11667 17085
rect 12894 17076 12900 17128
rect 12952 17116 12958 17128
rect 13446 17116 13452 17128
rect 12952 17088 13452 17116
rect 12952 17076 12958 17088
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 12802 17048 12808 17060
rect 12268 17020 12808 17048
rect 10870 16980 10876 16992
rect 10244 16952 10876 16980
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 12268 16980 12296 17020
rect 12802 17008 12808 17020
rect 12860 17048 12866 17060
rect 12860 17020 13400 17048
rect 12860 17008 12866 17020
rect 13372 16992 13400 17020
rect 11756 16952 12296 16980
rect 12621 16983 12679 16989
rect 11756 16940 11762 16952
rect 12621 16949 12633 16983
rect 12667 16980 12679 16983
rect 12710 16980 12716 16992
rect 12667 16952 12716 16980
rect 12667 16949 12679 16952
rect 12621 16943 12679 16949
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 13354 16940 13360 16992
rect 13412 16940 13418 16992
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 2498 16776 2504 16788
rect 1452 16748 2504 16776
rect 1452 16736 1458 16748
rect 2498 16736 2504 16748
rect 2556 16776 2562 16788
rect 2556 16748 2774 16776
rect 2556 16736 2562 16748
rect 2746 16640 2774 16748
rect 6730 16736 6736 16788
rect 6788 16776 6794 16788
rect 7098 16776 7104 16788
rect 6788 16748 7104 16776
rect 6788 16736 6794 16748
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 7745 16779 7803 16785
rect 7745 16745 7757 16779
rect 7791 16776 7803 16779
rect 8294 16776 8300 16788
rect 7791 16748 8300 16776
rect 7791 16745 7803 16748
rect 7745 16739 7803 16745
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 11790 16736 11796 16788
rect 11848 16736 11854 16788
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 14366 16776 14372 16788
rect 12584 16748 14372 16776
rect 12584 16736 12590 16748
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 8938 16668 8944 16720
rect 8996 16708 9002 16720
rect 10597 16711 10655 16717
rect 10597 16708 10609 16711
rect 8996 16680 10609 16708
rect 8996 16668 9002 16680
rect 10597 16677 10609 16680
rect 10643 16677 10655 16711
rect 10597 16671 10655 16677
rect 13725 16711 13783 16717
rect 13725 16677 13737 16711
rect 13771 16708 13783 16711
rect 13906 16708 13912 16720
rect 13771 16680 13912 16708
rect 13771 16677 13783 16680
rect 13725 16671 13783 16677
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 5994 16640 6000 16652
rect 2746 16612 6000 16640
rect 5994 16600 6000 16612
rect 6052 16640 6058 16652
rect 6730 16640 6736 16652
rect 6052 16612 6736 16640
rect 6052 16600 6058 16612
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10318 16640 10324 16652
rect 9999 16612 10324 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10870 16600 10876 16652
rect 10928 16600 10934 16652
rect 10990 16643 11048 16649
rect 10990 16609 11002 16643
rect 11036 16640 11048 16643
rect 11698 16640 11704 16652
rect 11036 16612 11704 16640
rect 11036 16609 11048 16612
rect 10990 16603 11048 16609
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 11790 16600 11796 16652
rect 11848 16640 11854 16652
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11848 16612 11897 16640
rect 11848 16600 11854 16612
rect 11885 16609 11897 16612
rect 11931 16640 11943 16643
rect 11974 16640 11980 16652
rect 11931 16612 11980 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 1394 16532 1400 16584
rect 1452 16532 1458 16584
rect 1671 16575 1729 16581
rect 1671 16541 1683 16575
rect 1717 16572 1729 16575
rect 1762 16572 1768 16584
rect 1717 16544 1768 16572
rect 1717 16541 1729 16544
rect 1671 16535 1729 16541
rect 1762 16532 1768 16544
rect 1820 16532 1826 16584
rect 7007 16575 7065 16581
rect 7007 16541 7019 16575
rect 7053 16572 7065 16575
rect 8662 16572 8668 16584
rect 7053 16544 8668 16572
rect 7053 16541 7065 16544
rect 7007 16535 7065 16541
rect 8662 16532 8668 16544
rect 8720 16572 8726 16584
rect 8846 16572 8852 16584
rect 8720 16544 8852 16572
rect 8720 16532 8726 16544
rect 8846 16532 8852 16544
rect 8904 16532 8910 16584
rect 10134 16532 10140 16584
rect 10192 16532 10198 16584
rect 11146 16532 11152 16584
rect 11204 16532 11210 16584
rect 12084 16572 12112 16603
rect 12526 16600 12532 16652
rect 12584 16600 12590 16652
rect 11900 16544 12112 16572
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 5718 16504 5724 16516
rect 3936 16476 5724 16504
rect 3936 16464 3942 16476
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 9582 16504 9588 16516
rect 6564 16476 9588 16504
rect 6564 16448 6592 16476
rect 9582 16464 9588 16476
rect 9640 16464 9646 16516
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 2409 16439 2467 16445
rect 2409 16436 2421 16439
rect 2004 16408 2421 16436
rect 2004 16396 2010 16408
rect 2409 16405 2421 16408
rect 2455 16405 2467 16439
rect 2409 16399 2467 16405
rect 6546 16396 6552 16448
rect 6604 16396 6610 16448
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 8478 16436 8484 16448
rect 7156 16408 8484 16436
rect 7156 16396 7162 16408
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 10152 16436 10180 16532
rect 11900 16436 11928 16544
rect 12802 16532 12808 16584
rect 12860 16532 12866 16584
rect 12894 16532 12900 16584
rect 12952 16581 12958 16584
rect 12952 16575 12980 16581
rect 12968 16541 12980 16575
rect 12952 16535 12980 16541
rect 12952 16532 12958 16535
rect 13078 16532 13084 16584
rect 13136 16532 13142 16584
rect 14274 16532 14280 16584
rect 14332 16532 14338 16584
rect 13722 16464 13728 16516
rect 13780 16504 13786 16516
rect 14461 16507 14519 16513
rect 14461 16504 14473 16507
rect 13780 16476 14473 16504
rect 13780 16464 13786 16476
rect 14461 16473 14473 16476
rect 14507 16473 14519 16507
rect 14461 16467 14519 16473
rect 10152 16408 11928 16436
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 12802 16436 12808 16448
rect 12492 16408 12808 16436
rect 12492 16396 12498 16408
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 6638 16192 6644 16244
rect 6696 16232 6702 16244
rect 7098 16232 7104 16244
rect 6696 16204 7104 16232
rect 6696 16192 6702 16204
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 11974 16232 11980 16244
rect 8772 16204 11980 16232
rect 7116 16164 7144 16192
rect 8202 16164 8208 16176
rect 7116 16136 8208 16164
rect 1655 16129 1713 16135
rect 1655 16095 1667 16129
rect 1701 16126 1713 16129
rect 1701 16096 1716 16126
rect 8202 16124 8208 16136
rect 8260 16164 8266 16176
rect 8260 16136 8616 16164
rect 8260 16124 8266 16136
rect 2038 16096 2044 16108
rect 1701 16095 2044 16096
rect 1655 16089 2044 16095
rect 1688 16068 2044 16089
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 7435 16099 7493 16105
rect 7435 16096 7447 16099
rect 6696 16068 7447 16096
rect 6696 16056 6702 16068
rect 7435 16065 7447 16068
rect 7481 16096 7493 16099
rect 7558 16096 7564 16108
rect 7481 16068 7564 16096
rect 7481 16065 7493 16068
rect 7435 16059 7493 16065
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8588 16105 8616 16136
rect 8772 16105 8800 16204
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 12526 16192 12532 16244
rect 12584 16192 12590 16244
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16201 14519 16235
rect 14461 16195 14519 16201
rect 10410 16124 10416 16176
rect 10468 16124 10474 16176
rect 14476 16164 14504 16195
rect 10980 16136 14504 16164
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 8573 16059 8631 16065
rect 8757 16099 8815 16105
rect 8757 16065 8769 16099
rect 8803 16065 8815 16099
rect 8757 16059 8815 16065
rect 8938 16056 8944 16108
rect 8996 16056 9002 16108
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 10980 16096 11008 16136
rect 10836 16068 11008 16096
rect 10836 16056 10842 16068
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11759 16099 11817 16105
rect 11759 16096 11771 16099
rect 11112 16068 11771 16096
rect 11112 16056 11118 16068
rect 11759 16065 11771 16068
rect 11805 16096 11817 16099
rect 13139 16099 13197 16105
rect 13139 16096 13151 16099
rect 11805 16068 13151 16096
rect 11805 16065 11817 16068
rect 11759 16059 11817 16065
rect 13139 16065 13151 16068
rect 13185 16065 13197 16099
rect 13139 16059 13197 16065
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16096 14335 16099
rect 15470 16096 15476 16108
rect 14323 16068 15476 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 15930 16096 15936 16108
rect 15804 16068 15936 16096
rect 15804 16056 15810 16068
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 1394 15988 1400 16040
rect 1452 15988 1458 16040
rect 6730 15988 6736 16040
rect 6788 16028 6794 16040
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 6788 16000 7205 16028
rect 6788 15988 6794 16000
rect 7193 15997 7205 16000
rect 7239 15997 7251 16031
rect 8956 16028 8984 16056
rect 9493 16031 9551 16037
rect 9493 16028 9505 16031
rect 7193 15991 7251 15997
rect 8128 16000 9505 16028
rect 6914 15920 6920 15972
rect 6972 15920 6978 15972
rect 2406 15852 2412 15904
rect 2464 15852 2470 15904
rect 6932 15892 6960 15920
rect 8128 15892 8156 16000
rect 9493 15997 9505 16000
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 9582 15988 9588 16040
rect 9640 16037 9646 16040
rect 9640 16031 9668 16037
rect 9656 15997 9668 16031
rect 9640 15991 9668 15997
rect 9640 15988 9646 15991
rect 9766 15988 9772 16040
rect 9824 15988 9830 16040
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 11146 16028 11152 16040
rect 10468 16000 11152 16028
rect 10468 15988 10474 16000
rect 11146 15988 11152 16000
rect 11204 16028 11210 16040
rect 11514 16028 11520 16040
rect 11204 16000 11520 16028
rect 11204 15988 11210 16000
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 12802 16028 12808 16040
rect 12400 16000 12808 16028
rect 12400 15988 12406 16000
rect 12802 15988 12808 16000
rect 12860 16028 12866 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12860 16000 12909 16028
rect 12860 15988 12866 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 8205 15963 8263 15969
rect 8205 15929 8217 15963
rect 8251 15960 8263 15963
rect 9217 15963 9275 15969
rect 9217 15960 9229 15963
rect 8251 15932 9229 15960
rect 8251 15929 8263 15932
rect 8205 15923 8263 15929
rect 9217 15929 9229 15932
rect 9263 15929 9275 15963
rect 9217 15923 9275 15929
rect 12434 15920 12440 15972
rect 12492 15960 12498 15972
rect 12492 15932 12940 15960
rect 12492 15920 12498 15932
rect 6932 15864 8156 15892
rect 9122 15852 9128 15904
rect 9180 15892 9186 15904
rect 11146 15892 11152 15904
rect 9180 15864 11152 15892
rect 9180 15852 9186 15864
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11606 15852 11612 15904
rect 11664 15892 11670 15904
rect 12802 15892 12808 15904
rect 11664 15864 12808 15892
rect 11664 15852 11670 15864
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 12912 15892 12940 15932
rect 13556 15892 13584 16056
rect 12912 15864 13584 15892
rect 13906 15852 13912 15904
rect 13964 15852 13970 15904
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 5350 15688 5356 15700
rect 1627 15660 5356 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 5552 15660 9904 15688
rect 2314 15580 2320 15632
rect 2372 15620 2378 15632
rect 5552 15620 5580 15660
rect 2372 15592 5580 15620
rect 2372 15580 2378 15592
rect 6362 15580 6368 15632
rect 6420 15620 6426 15632
rect 6914 15620 6920 15632
rect 6420 15592 6920 15620
rect 6420 15580 6426 15592
rect 6914 15580 6920 15592
rect 6972 15580 6978 15632
rect 9876 15620 9904 15660
rect 9950 15648 9956 15700
rect 10008 15648 10014 15700
rect 11054 15688 11060 15700
rect 10428 15660 11060 15688
rect 10428 15620 10456 15660
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 13906 15688 13912 15700
rect 11204 15660 12296 15688
rect 11204 15648 11210 15660
rect 11977 15623 12035 15629
rect 11977 15620 11989 15623
rect 9876 15592 10456 15620
rect 10980 15592 11989 15620
rect 8570 15512 8576 15564
rect 8628 15552 8634 15564
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8628 15524 8953 15552
rect 8628 15512 8634 15524
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 750 15444 756 15496
rect 808 15484 814 15496
rect 1489 15487 1547 15493
rect 1489 15484 1501 15487
rect 808 15456 1501 15484
rect 808 15444 814 15456
rect 1489 15453 1501 15456
rect 1535 15453 1547 15487
rect 1489 15447 1547 15453
rect 1578 15444 1584 15496
rect 1636 15444 1642 15496
rect 1946 15444 1952 15496
rect 2004 15444 2010 15496
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 5132 15456 5457 15484
rect 5132 15444 5138 15456
rect 5445 15453 5457 15456
rect 5491 15453 5503 15487
rect 9214 15484 9220 15496
rect 5703 15477 5761 15483
rect 5703 15474 5715 15477
rect 5445 15447 5503 15453
rect 5644 15446 5715 15474
rect 1596 15416 1624 15444
rect 5644 15416 5672 15446
rect 5703 15443 5715 15446
rect 5749 15443 5761 15477
rect 9175 15456 9220 15484
rect 9214 15444 9220 15456
rect 9272 15444 9278 15496
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 9824 15456 10333 15484
rect 9824 15444 9830 15456
rect 10321 15453 10333 15456
rect 10367 15484 10379 15487
rect 10980 15484 11008 15592
rect 11977 15589 11989 15592
rect 12023 15589 12035 15623
rect 11977 15583 12035 15589
rect 12268 15561 12296 15660
rect 12728 15660 13912 15688
rect 12728 15629 12756 15660
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 14366 15648 14372 15700
rect 14424 15648 14430 15700
rect 12713 15623 12771 15629
rect 12713 15589 12725 15623
rect 12759 15589 12771 15623
rect 12713 15583 12771 15589
rect 12253 15555 12311 15561
rect 11808 15524 12204 15552
rect 11808 15493 11836 15524
rect 10367 15456 10456 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 5703 15437 5761 15443
rect 10428 15428 10456 15456
rect 10579 15457 10637 15463
rect 8294 15416 8300 15428
rect 1596 15388 5672 15416
rect 6380 15388 8300 15416
rect 1762 15308 1768 15360
rect 1820 15308 1826 15360
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 6380 15348 6408 15388
rect 8294 15376 8300 15388
rect 8352 15376 8358 15428
rect 10410 15376 10416 15428
rect 10468 15376 10474 15428
rect 10579 15423 10591 15457
rect 10625 15454 10637 15457
rect 10704 15456 11008 15484
rect 11793 15487 11851 15493
rect 10625 15423 10640 15454
rect 10579 15417 10640 15423
rect 5408 15320 6408 15348
rect 5408 15308 5414 15320
rect 6454 15308 6460 15360
rect 6512 15308 6518 15360
rect 8754 15308 8760 15360
rect 8812 15348 8818 15360
rect 9214 15348 9220 15360
rect 8812 15320 9220 15348
rect 8812 15308 8818 15320
rect 9214 15308 9220 15320
rect 9272 15348 9278 15360
rect 10612 15348 10640 15417
rect 10704 15416 10732 15456
rect 11793 15453 11805 15487
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15453 12127 15487
rect 12176 15484 12204 15524
rect 12253 15521 12265 15555
rect 12299 15521 12311 15555
rect 14090 15552 14096 15564
rect 12253 15515 12311 15521
rect 12406 15524 14096 15552
rect 12406 15484 12434 15524
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 12176 15456 12434 15484
rect 12069 15447 12127 15453
rect 10778 15416 10784 15428
rect 10704 15388 10784 15416
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 12084 15416 12112 15447
rect 12986 15444 12992 15496
rect 13044 15444 13050 15496
rect 13078 15444 13084 15496
rect 13136 15493 13142 15496
rect 13136 15487 13164 15493
rect 13152 15453 13164 15487
rect 13136 15447 13164 15453
rect 13136 15444 13142 15447
rect 13262 15444 13268 15496
rect 13320 15444 13326 15496
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 14550 15484 14556 15496
rect 14323 15456 14556 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 10888 15388 12112 15416
rect 13909 15419 13967 15425
rect 9272 15320 10640 15348
rect 9272 15308 9278 15320
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 10888 15348 10916 15388
rect 13909 15385 13921 15419
rect 13955 15416 13967 15419
rect 15764 15416 15792 15444
rect 13955 15388 15792 15416
rect 13955 15385 13967 15388
rect 13909 15379 13967 15385
rect 10744 15320 10916 15348
rect 11333 15351 11391 15357
rect 10744 15308 10750 15320
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 11606 15348 11612 15360
rect 11379 15320 11612 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 13078 15348 13084 15360
rect 12032 15320 13084 15348
rect 12032 15308 12038 15320
rect 13078 15308 13084 15320
rect 13136 15308 13142 15360
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 2406 15104 2412 15156
rect 2464 15104 2470 15156
rect 6546 15104 6552 15156
rect 6604 15104 6610 15156
rect 6730 15104 6736 15156
rect 6788 15144 6794 15156
rect 7653 15147 7711 15153
rect 7653 15144 7665 15147
rect 6788 15116 7665 15144
rect 6788 15104 6794 15116
rect 7653 15113 7665 15116
rect 7699 15113 7711 15147
rect 7653 15107 7711 15113
rect 7837 15147 7895 15153
rect 7837 15113 7849 15147
rect 7883 15144 7895 15147
rect 8202 15144 8208 15156
rect 7883 15116 8208 15144
rect 7883 15113 7895 15116
rect 7837 15107 7895 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8352 15116 9674 15144
rect 8352 15104 8358 15116
rect 1489 15079 1547 15085
rect 1489 15045 1501 15079
rect 1535 15076 1547 15079
rect 1762 15076 1768 15088
rect 1535 15048 1768 15076
rect 1535 15045 1547 15048
rect 1489 15039 1547 15045
rect 1762 15036 1768 15048
rect 1820 15036 1826 15088
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 15008 2191 15011
rect 2424 15008 2452 15104
rect 6362 15036 6368 15088
rect 6420 15076 6426 15088
rect 6825 15079 6883 15085
rect 6825 15076 6837 15079
rect 6420 15048 6837 15076
rect 6420 15036 6426 15048
rect 6825 15045 6837 15048
rect 6871 15045 6883 15079
rect 9646 15076 9674 15116
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12676 15116 12817 15144
rect 12676 15104 12682 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 14001 15147 14059 15153
rect 14001 15144 14013 15147
rect 13320 15116 14013 15144
rect 13320 15104 13326 15116
rect 14001 15113 14013 15116
rect 14047 15113 14059 15147
rect 14001 15107 14059 15113
rect 9646 15048 11744 15076
rect 6825 15039 6883 15045
rect 2179 14980 2452 15008
rect 2179 14977 2191 14980
rect 2133 14971 2191 14977
rect 6914 14968 6920 15020
rect 6972 14968 6978 15020
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 7156 14980 7297 15008
rect 7156 14968 7162 14980
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7285 14971 7343 14977
rect 9692 15008 9904 15018
rect 10011 15011 10069 15017
rect 10011 15008 10023 15011
rect 9692 14990 10023 15008
rect 6454 14900 6460 14952
rect 6512 14900 6518 14952
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 9692 14940 9720 14990
rect 9876 14980 10023 14990
rect 10011 14977 10023 14980
rect 10057 14977 10069 15011
rect 10011 14971 10069 14977
rect 8628 14912 9720 14940
rect 8628 14900 8634 14912
rect 9766 14900 9772 14952
rect 9824 14900 9830 14952
rect 10778 14940 10784 14952
rect 10704 14912 10784 14940
rect 8386 14832 8392 14884
rect 8444 14872 8450 14884
rect 9030 14872 9036 14884
rect 8444 14844 9036 14872
rect 8444 14832 8450 14844
rect 9030 14832 9036 14844
rect 9088 14832 9094 14884
rect 842 14764 848 14816
rect 900 14804 906 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 900 14776 1593 14804
rect 900 14764 906 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 1946 14764 1952 14816
rect 2004 14764 2010 14816
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 10226 14804 10232 14816
rect 10100 14776 10232 14804
rect 10100 14764 10106 14776
rect 10226 14764 10232 14776
rect 10284 14804 10290 14816
rect 10704 14804 10732 14912
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 10284 14776 10732 14804
rect 10284 14764 10290 14776
rect 10778 14764 10784 14816
rect 10836 14764 10842 14816
rect 11716 14804 11744 15048
rect 12066 15036 12072 15088
rect 12124 15076 12130 15088
rect 12713 15079 12771 15085
rect 12124 15048 12664 15076
rect 12124 15036 12130 15048
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 15008 11851 15011
rect 11974 15008 11980 15020
rect 11839 14980 11980 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12636 15008 12664 15048
rect 12713 15045 12725 15079
rect 12759 15076 12771 15079
rect 14182 15076 14188 15088
rect 12759 15048 14188 15076
rect 12759 15045 12771 15048
rect 12713 15039 12771 15045
rect 14182 15036 14188 15048
rect 14240 15036 14246 15088
rect 13231 15011 13289 15017
rect 13231 15008 13243 15011
rect 12636 14980 13243 15008
rect 13231 14977 13243 14980
rect 13277 14977 13289 15011
rect 13231 14971 13289 14977
rect 12526 14940 12532 14952
rect 11992 14912 12532 14940
rect 11992 14884 12020 14912
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 12989 14943 13047 14949
rect 12989 14940 13001 14943
rect 12768 14912 13001 14940
rect 12768 14900 12774 14912
rect 12989 14909 13001 14912
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 11974 14832 11980 14884
rect 12032 14832 12038 14884
rect 12066 14832 12072 14884
rect 12124 14872 12130 14884
rect 12434 14872 12440 14884
rect 12124 14844 12440 14872
rect 12124 14832 12130 14844
rect 12434 14832 12440 14844
rect 12492 14832 12498 14884
rect 14550 14804 14556 14816
rect 11716 14776 14556 14804
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 6825 14603 6883 14609
rect 5828 14572 6776 14600
rect 3786 14492 3792 14544
rect 3844 14532 3850 14544
rect 5626 14532 5632 14544
rect 3844 14504 5632 14532
rect 3844 14492 3850 14504
rect 5626 14492 5632 14504
rect 5684 14492 5690 14544
rect 5074 14424 5080 14476
rect 5132 14464 5138 14476
rect 5534 14464 5540 14476
rect 5132 14436 5540 14464
rect 5132 14424 5138 14436
rect 5534 14424 5540 14436
rect 5592 14464 5598 14476
rect 5828 14473 5856 14572
rect 5813 14467 5871 14473
rect 5813 14464 5825 14467
rect 5592 14436 5825 14464
rect 5592 14424 5598 14436
rect 5813 14433 5825 14436
rect 5859 14433 5871 14467
rect 5813 14427 5871 14433
rect 1394 14356 1400 14408
rect 1452 14356 1458 14408
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 6055 14399 6113 14405
rect 6055 14396 6067 14399
rect 1728 14368 4476 14396
rect 1728 14356 1734 14368
rect 1210 14288 1216 14340
rect 1268 14328 1274 14340
rect 4448 14328 4476 14368
rect 5920 14368 6067 14396
rect 5920 14328 5948 14368
rect 6055 14365 6067 14368
rect 6101 14365 6113 14399
rect 6748 14396 6776 14572
rect 6825 14569 6837 14603
rect 6871 14600 6883 14603
rect 6914 14600 6920 14612
rect 6871 14572 6920 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 7208 14572 8984 14600
rect 7208 14544 7236 14572
rect 7190 14492 7196 14544
rect 7248 14492 7254 14544
rect 8956 14464 8984 14572
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 9398 14600 9404 14612
rect 9180 14572 9404 14600
rect 9180 14560 9186 14572
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 10836 14572 11100 14600
rect 10836 14560 10842 14572
rect 9582 14492 9588 14544
rect 9640 14532 9646 14544
rect 11072 14541 11100 14572
rect 11514 14560 11520 14612
rect 11572 14600 11578 14612
rect 11790 14600 11796 14612
rect 11572 14572 11796 14600
rect 11572 14560 11578 14572
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 12158 14560 12164 14612
rect 12216 14600 12222 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 12216 14572 12265 14600
rect 12216 14560 12222 14572
rect 12253 14569 12265 14572
rect 12299 14569 12311 14603
rect 12253 14563 12311 14569
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 14369 14603 14427 14609
rect 14369 14600 14381 14603
rect 13504 14572 14381 14600
rect 13504 14560 13510 14572
rect 14369 14569 14381 14572
rect 14415 14569 14427 14603
rect 14369 14563 14427 14569
rect 11057 14535 11115 14541
rect 9640 14504 10824 14532
rect 9640 14492 9646 14504
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 8956 14436 10425 14464
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 7193 14399 7251 14405
rect 7193 14396 7205 14399
rect 6748 14368 7205 14396
rect 6055 14359 6113 14365
rect 7193 14365 7205 14368
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 7467 14399 7525 14405
rect 7467 14365 7479 14399
rect 7513 14396 7525 14399
rect 7513 14368 7880 14396
rect 7513 14365 7525 14368
rect 7467 14359 7525 14365
rect 1268 14300 2774 14328
rect 4448 14300 5948 14328
rect 1268 14288 1274 14300
rect 2406 14220 2412 14272
rect 2464 14220 2470 14272
rect 2746 14260 2774 14300
rect 7098 14260 7104 14272
rect 2746 14232 7104 14260
rect 7098 14220 7104 14232
rect 7156 14260 7162 14272
rect 7852 14260 7880 14368
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 9766 14396 9772 14408
rect 8904 14368 9772 14396
rect 8904 14356 8910 14368
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 10428 14396 10456 14427
rect 10502 14424 10508 14476
rect 10560 14464 10566 14476
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 10560 14436 10609 14464
rect 10560 14424 10566 14436
rect 10597 14433 10609 14436
rect 10643 14464 10655 14467
rect 10686 14464 10692 14476
rect 10643 14436 10692 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 10796 14464 10824 14504
rect 11057 14501 11069 14535
rect 11103 14501 11115 14535
rect 11057 14495 11115 14501
rect 11146 14464 11152 14476
rect 10796 14436 11152 14464
rect 11146 14424 11152 14436
rect 11204 14464 11210 14476
rect 11450 14467 11508 14473
rect 11450 14464 11462 14467
rect 11204 14436 11462 14464
rect 11204 14424 11210 14436
rect 11450 14433 11462 14436
rect 11496 14433 11508 14467
rect 11450 14427 11508 14433
rect 11606 14424 11612 14476
rect 11664 14424 11670 14476
rect 11974 14424 11980 14476
rect 12032 14464 12038 14476
rect 12032 14436 12204 14464
rect 12032 14424 12038 14436
rect 10778 14396 10784 14408
rect 10428 14368 10784 14396
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11330 14356 11336 14408
rect 11388 14356 11394 14408
rect 12176 14396 12204 14436
rect 12618 14424 12624 14476
rect 12676 14424 12682 14476
rect 12342 14396 12348 14408
rect 12176 14368 12348 14396
rect 12342 14356 12348 14368
rect 12400 14396 12406 14408
rect 12863 14399 12921 14405
rect 12863 14396 12875 14399
rect 12400 14368 12875 14396
rect 12400 14356 12406 14368
rect 12863 14365 12875 14368
rect 12909 14365 12921 14399
rect 12863 14359 12921 14365
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 13780 14368 14289 14396
rect 13780 14356 13786 14368
rect 14277 14365 14289 14368
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 8294 14288 8300 14340
rect 8352 14328 8358 14340
rect 8478 14328 8484 14340
rect 8352 14300 8484 14328
rect 8352 14288 8358 14300
rect 8478 14288 8484 14300
rect 8536 14328 8542 14340
rect 9582 14328 9588 14340
rect 8536 14300 9588 14328
rect 8536 14288 8542 14300
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 13372 14300 14412 14328
rect 7156 14232 7880 14260
rect 7156 14220 7162 14232
rect 8202 14220 8208 14272
rect 8260 14220 8266 14272
rect 8846 14220 8852 14272
rect 8904 14260 8910 14272
rect 11330 14260 11336 14272
rect 8904 14232 11336 14260
rect 8904 14220 8910 14232
rect 11330 14220 11336 14232
rect 11388 14260 11394 14272
rect 13372 14260 13400 14300
rect 14384 14272 14412 14300
rect 11388 14232 13400 14260
rect 13633 14263 13691 14269
rect 11388 14220 11394 14232
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 13814 14260 13820 14272
rect 13679 14232 13820 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 14366 14220 14372 14272
rect 14424 14220 14430 14272
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 842 14016 848 14068
rect 900 14056 906 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 900 14028 1593 14056
rect 900 14016 906 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 1581 14019 1639 14025
rect 1946 14016 1952 14068
rect 2004 14016 2010 14068
rect 2406 14016 2412 14068
rect 2464 14016 2470 14068
rect 7098 14016 7104 14068
rect 7156 14016 7162 14068
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 8757 14059 8815 14065
rect 7892 14028 8708 14056
rect 7892 14016 7898 14028
rect 1489 13991 1547 13997
rect 1489 13957 1501 13991
rect 1535 13988 1547 13991
rect 1964 13988 1992 14016
rect 1535 13960 1992 13988
rect 1535 13957 1547 13960
rect 1489 13951 1547 13957
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2424 13920 2452 14016
rect 2179 13892 2452 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 5810 13880 5816 13932
rect 5868 13880 5874 13932
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13920 6975 13923
rect 7116 13920 7144 14016
rect 8680 13988 8708 14028
rect 8757 14025 8769 14059
rect 8803 14056 8815 14059
rect 9306 14056 9312 14068
rect 8803 14028 9312 14056
rect 8803 14025 8815 14028
rect 8757 14019 8815 14025
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 10321 14059 10379 14065
rect 10321 14025 10333 14059
rect 10367 14056 10379 14059
rect 12066 14056 12072 14068
rect 10367 14028 12072 14056
rect 10367 14025 10379 14028
rect 10321 14019 10379 14025
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 12250 14016 12256 14068
rect 12308 14056 12314 14068
rect 13630 14056 13636 14068
rect 12308 14028 13636 14056
rect 12308 14016 12314 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 14461 14059 14519 14065
rect 14461 14025 14473 14059
rect 14507 14056 14519 14059
rect 15194 14056 15200 14068
rect 14507 14028 15200 14056
rect 14507 14025 14519 14028
rect 14461 14019 14519 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 8846 13988 8852 14000
rect 8680 13960 8852 13988
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 9030 13948 9036 14000
rect 9088 13948 9094 14000
rect 10042 13988 10048 14000
rect 9324 13960 10048 13988
rect 6963 13892 7144 13920
rect 6963 13889 6975 13892
rect 6917 13883 6975 13889
rect 8110 13880 8116 13932
rect 8168 13880 8174 13932
rect 9324 13929 9352 13960
rect 10042 13948 10048 13960
rect 10100 13948 10106 14000
rect 10137 13991 10195 13997
rect 10137 13957 10149 13991
rect 10183 13988 10195 13991
rect 11054 13988 11060 14000
rect 10183 13960 11060 13988
rect 10183 13957 10195 13960
rect 10137 13951 10195 13957
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 11698 13988 11704 14000
rect 11532 13960 11704 13988
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13889 9367 13923
rect 9309 13883 9367 13889
rect 9398 13880 9404 13932
rect 9456 13880 9462 13932
rect 9766 13880 9772 13932
rect 9824 13920 9830 13932
rect 10226 13920 10232 13932
rect 9824 13892 10232 13920
rect 9824 13880 9830 13892
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 11532 13929 11560 13960
rect 11698 13948 11704 13960
rect 11756 13988 11762 14000
rect 11974 13988 11980 14000
rect 11756 13960 11980 13988
rect 11756 13948 11762 13960
rect 11974 13948 11980 13960
rect 12032 13948 12038 14000
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13889 11575 13923
rect 11790 13920 11796 13932
rect 11751 13892 11796 13920
rect 11517 13883 11575 13889
rect 11790 13880 11796 13892
rect 11848 13920 11854 13932
rect 13139 13923 13197 13929
rect 13139 13920 13151 13923
rect 11848 13892 13151 13920
rect 11848 13880 11854 13892
rect 13139 13889 13151 13892
rect 13185 13889 13197 13923
rect 13139 13883 13197 13889
rect 14274 13880 14280 13932
rect 14332 13880 14338 13932
rect 566 13812 572 13864
rect 624 13852 630 13864
rect 4246 13852 4252 13864
rect 624 13824 4252 13852
rect 624 13812 630 13824
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 5828 13852 5856 13880
rect 7101 13855 7159 13861
rect 5828 13824 7052 13852
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 5810 13784 5816 13796
rect 5500 13756 5816 13784
rect 5500 13744 5506 13756
rect 5810 13744 5816 13756
rect 5868 13744 5874 13796
rect 7024 13784 7052 13824
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7190 13852 7196 13864
rect 7147 13824 7196 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 7834 13852 7840 13864
rect 7484 13824 7840 13852
rect 7484 13784 7512 13824
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 7975 13855 8033 13861
rect 7975 13821 7987 13855
rect 8021 13852 8033 13855
rect 8294 13852 8300 13864
rect 8021 13824 8300 13852
rect 8021 13821 8033 13824
rect 7975 13815 8033 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8536 13824 8878 13852
rect 8536 13812 8542 13824
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12676 13824 12909 13852
rect 12676 13812 12682 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 7024 13756 7512 13784
rect 7558 13744 7564 13796
rect 7616 13744 7622 13796
rect 12636 13784 12664 13812
rect 12176 13756 12664 13784
rect 1946 13676 1952 13728
rect 2004 13676 2010 13728
rect 7374 13676 7380 13728
rect 7432 13716 7438 13728
rect 9030 13716 9036 13728
rect 7432 13688 9036 13716
rect 7432 13676 7438 13688
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 12176 13716 12204 13756
rect 13998 13744 14004 13796
rect 14056 13784 14062 13796
rect 14274 13784 14280 13796
rect 14056 13756 14280 13784
rect 14056 13744 14062 13756
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 10744 13688 12204 13716
rect 10744 13676 10750 13688
rect 12526 13676 12532 13728
rect 12584 13676 12590 13728
rect 13262 13676 13268 13728
rect 13320 13716 13326 13728
rect 13909 13719 13967 13725
rect 13909 13716 13921 13719
rect 13320 13688 13921 13716
rect 13320 13676 13326 13688
rect 13909 13685 13921 13688
rect 13955 13685 13967 13719
rect 13909 13679 13967 13685
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 7101 13515 7159 13521
rect 6104 13484 7052 13512
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 6104 13385 6132 13484
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5592 13348 6101 13376
rect 5592 13336 5598 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 7024 13376 7052 13484
rect 7101 13481 7113 13515
rect 7147 13512 7159 13515
rect 7558 13512 7564 13524
rect 7147 13484 7564 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 8478 13472 8484 13524
rect 8536 13472 8542 13524
rect 9398 13472 9404 13524
rect 9456 13512 9462 13524
rect 9953 13515 10011 13521
rect 9953 13512 9965 13515
rect 9456 13484 9965 13512
rect 9456 13472 9462 13484
rect 9953 13481 9965 13484
rect 9999 13481 10011 13515
rect 12526 13512 12532 13524
rect 9953 13475 10011 13481
rect 12176 13484 12532 13512
rect 12176 13453 12204 13484
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 12952 13484 13369 13512
rect 12952 13472 12958 13484
rect 13357 13481 13369 13484
rect 13403 13481 13415 13515
rect 13357 13475 13415 13481
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 14274 13512 14280 13524
rect 13955 13484 14280 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 14366 13472 14372 13524
rect 14424 13472 14430 13524
rect 12161 13447 12219 13453
rect 12161 13413 12173 13447
rect 12207 13413 12219 13447
rect 13446 13444 13452 13456
rect 12161 13407 12219 13413
rect 13372 13416 13452 13444
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7024 13348 7481 13376
rect 6089 13339 6147 13345
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 1489 13311 1547 13317
rect 1489 13277 1501 13311
rect 1535 13308 1547 13311
rect 1946 13308 1952 13320
rect 1535 13280 1952 13308
rect 1535 13277 1547 13280
rect 1489 13271 1547 13277
rect 1946 13268 1952 13280
rect 2004 13268 2010 13320
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 5868 13281 6408 13308
rect 5868 13280 6359 13281
rect 5868 13268 5874 13280
rect 6347 13247 6359 13280
rect 6393 13250 6408 13281
rect 6393 13247 6405 13250
rect 6347 13241 6405 13247
rect 842 13132 848 13184
rect 900 13172 906 13184
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 900 13144 1593 13172
rect 900 13132 906 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 7484 13172 7512 13339
rect 10042 13336 10048 13388
rect 10100 13376 10106 13388
rect 10318 13376 10324 13388
rect 10100 13348 10324 13376
rect 10100 13336 10106 13348
rect 10318 13336 10324 13348
rect 10376 13376 10382 13388
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 10376 13348 11713 13376
rect 10376 13336 10382 13348
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 11882 13336 11888 13388
rect 11940 13336 11946 13388
rect 12250 13336 12256 13388
rect 12308 13376 12314 13388
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 12308 13348 12449 13376
rect 12308 13336 12314 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12575 13379 12633 13385
rect 12575 13345 12587 13379
rect 12621 13376 12633 13379
rect 13372 13376 13400 13416
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 14642 13376 14648 13388
rect 12621 13348 13400 13376
rect 13464 13348 14648 13376
rect 12621 13345 12633 13348
rect 12575 13339 12633 13345
rect 7743 13311 7801 13317
rect 7743 13277 7755 13311
rect 7789 13308 7801 13311
rect 7789 13280 8248 13308
rect 7789 13277 7801 13280
rect 7743 13271 7801 13277
rect 8220 13252 8248 13280
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 8846 13308 8852 13320
rect 8628 13280 8852 13308
rect 8628 13268 8634 13280
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9215 13311 9273 13317
rect 9215 13277 9227 13311
rect 9261 13308 9273 13311
rect 9261 13280 9444 13308
rect 9261 13277 9273 13280
rect 9215 13271 9273 13277
rect 8202 13200 8208 13252
rect 8260 13200 8266 13252
rect 8956 13172 8984 13271
rect 9416 13252 9444 13280
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11204 13280 11529 13308
rect 11204 13268 11210 13280
rect 11517 13277 11529 13280
rect 11563 13308 11575 13311
rect 11900 13308 11928 13336
rect 11563 13280 11928 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 13464 13317 13492 13348
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 13722 13268 13728 13320
rect 13780 13268 13786 13320
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 15654 13308 15660 13320
rect 14323 13280 15660 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 9398 13200 9404 13252
rect 9456 13200 9462 13252
rect 13188 13212 13676 13240
rect 9858 13172 9864 13184
rect 7484 13144 9864 13172
rect 1581 13135 1639 13141
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 13188 13172 13216 13212
rect 13648 13181 13676 13212
rect 11296 13144 13216 13172
rect 13633 13175 13691 13181
rect 11296 13132 11302 13144
rect 13633 13141 13645 13175
rect 13679 13141 13691 13175
rect 13633 13135 13691 13141
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 15838 13172 15844 13184
rect 13780 13144 15844 13172
rect 13780 13132 13786 13144
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 1578 12928 1584 12980
rect 1636 12968 1642 12980
rect 1636 12940 1716 12968
rect 1636 12928 1642 12940
rect 1688 12851 1716 12940
rect 4706 12928 4712 12980
rect 4764 12968 4770 12980
rect 8570 12968 8576 12980
rect 4764 12940 8576 12968
rect 4764 12928 4770 12940
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11756 12940 11989 12968
rect 11756 12928 11762 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 15194 12968 15200 12980
rect 11977 12931 12035 12937
rect 12360 12940 15200 12968
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 7156 12872 9674 12900
rect 7156 12860 7162 12872
rect 1671 12845 1729 12851
rect 1671 12811 1683 12845
rect 1717 12811 1729 12845
rect 1671 12805 1729 12811
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 9398 12832 9404 12844
rect 6880 12804 9404 12832
rect 6880 12792 6886 12804
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 1394 12724 1400 12776
rect 1452 12724 1458 12776
rect 2406 12588 2412 12640
rect 2464 12588 2470 12640
rect 9646 12628 9674 12872
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 10778 12832 10784 12844
rect 10100 12804 10784 12832
rect 10100 12792 10106 12804
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 11054 12792 11060 12844
rect 11112 12792 11118 12844
rect 11790 12792 11796 12844
rect 11848 12792 11854 12844
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 12250 12832 12256 12844
rect 12115 12804 12256 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 12360 12841 12388 12940
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 12345 12835 12403 12841
rect 12345 12801 12357 12835
rect 12391 12801 12403 12835
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12345 12795 12403 12801
rect 12452 12804 12817 12832
rect 11072 12764 11100 12792
rect 12158 12764 12164 12776
rect 11072 12736 12164 12764
rect 12158 12724 12164 12736
rect 12216 12764 12222 12776
rect 12452 12764 12480 12804
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 12805 12795 12863 12801
rect 13538 12792 13544 12844
rect 13596 12792 13602 12844
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 12216 12736 12480 12764
rect 12216 12724 12222 12736
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 12584 12736 12633 12764
rect 12584 12724 12590 12736
rect 12621 12733 12633 12736
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 13630 12724 13636 12776
rect 13688 12773 13694 12776
rect 13688 12767 13716 12773
rect 13704 12733 13716 12767
rect 13688 12727 13716 12733
rect 13688 12724 13694 12727
rect 13262 12656 13268 12708
rect 13320 12656 13326 12708
rect 14458 12656 14464 12708
rect 14516 12656 14522 12708
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 9646 12600 12265 12628
rect 12253 12597 12265 12600
rect 12299 12597 12311 12631
rect 12253 12591 12311 12597
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12529 12631 12587 12637
rect 12529 12628 12541 12631
rect 12492 12600 12541 12628
rect 12492 12588 12498 12600
rect 12529 12597 12541 12600
rect 12575 12597 12587 12631
rect 12529 12591 12587 12597
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 842 12384 848 12436
rect 900 12424 906 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 900 12396 1593 12424
rect 900 12384 906 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 10686 12424 10692 12436
rect 9916 12396 10692 12424
rect 9916 12384 9922 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11882 12424 11888 12436
rect 11440 12396 11888 12424
rect 8754 12316 8760 12368
rect 8812 12356 8818 12368
rect 10410 12356 10416 12368
rect 8812 12328 10416 12356
rect 8812 12316 8818 12328
rect 10410 12316 10416 12328
rect 10468 12356 10474 12368
rect 10962 12356 10968 12368
rect 10468 12328 10968 12356
rect 10468 12316 10474 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5902 12288 5908 12300
rect 4948 12260 5908 12288
rect 4948 12248 4954 12260
rect 5902 12248 5908 12260
rect 5960 12288 5966 12300
rect 6549 12291 6607 12297
rect 6549 12288 6561 12291
rect 5960 12260 6561 12288
rect 5960 12248 5966 12260
rect 6549 12257 6561 12260
rect 6595 12257 6607 12291
rect 6549 12251 6607 12257
rect 10226 12248 10232 12300
rect 10284 12288 10290 12300
rect 10686 12288 10692 12300
rect 10284 12260 10692 12288
rect 10284 12248 10290 12260
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 11440 12297 11468 12396
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 12437 12427 12495 12433
rect 12437 12393 12449 12427
rect 12483 12424 12495 12427
rect 12710 12424 12716 12436
rect 12483 12396 12716 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 13906 12424 13912 12436
rect 13504 12396 13912 12424
rect 13504 12384 13510 12396
rect 13906 12384 13912 12396
rect 13964 12424 13970 12436
rect 15930 12424 15936 12436
rect 13964 12396 15936 12424
rect 13964 12384 13970 12396
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 14274 12316 14280 12368
rect 14332 12316 14338 12368
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 12805 12291 12863 12297
rect 12805 12257 12817 12291
rect 12851 12288 12863 12291
rect 14292 12288 14320 12316
rect 12851 12260 14320 12288
rect 12851 12257 12863 12260
rect 12805 12251 12863 12257
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2406 12220 2412 12232
rect 2179 12192 2412 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 6791 12223 6849 12229
rect 6791 12220 6803 12223
rect 6656 12192 6803 12220
rect 6656 12164 6684 12192
rect 6791 12189 6803 12192
rect 6837 12189 6849 12223
rect 6791 12183 6849 12189
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10594 12220 10600 12232
rect 9824 12192 10600 12220
rect 9824 12180 9830 12192
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 11699 12223 11757 12229
rect 11699 12189 11711 12223
rect 11745 12220 11757 12223
rect 12342 12220 12348 12232
rect 11745 12192 12348 12220
rect 11745 12189 11757 12192
rect 11699 12183 11757 12189
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13262 12220 13268 12232
rect 13127 12192 13268 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13262 12180 13268 12192
rect 13320 12220 13326 12232
rect 13446 12220 13452 12232
rect 13320 12192 13452 12220
rect 13320 12180 13326 12192
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 14182 12220 14188 12232
rect 13771 12192 14188 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 15470 12220 15476 12232
rect 14323 12192 15476 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 1489 12155 1547 12161
rect 1489 12121 1501 12155
rect 1535 12152 1547 12155
rect 1535 12124 1992 12152
rect 1535 12121 1547 12124
rect 1489 12115 1547 12121
rect 1964 12093 1992 12124
rect 6638 12112 6644 12164
rect 6696 12112 6702 12164
rect 9122 12112 9128 12164
rect 9180 12152 9186 12164
rect 9180 12124 14504 12152
rect 9180 12112 9186 12124
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12053 2007 12087
rect 1949 12047 2007 12053
rect 7558 12044 7564 12096
rect 7616 12044 7622 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 10318 12084 10324 12096
rect 9272 12056 10324 12084
rect 9272 12044 9278 12056
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 13814 12084 13820 12096
rect 11848 12056 13820 12084
rect 11848 12044 11854 12056
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 14476 12093 14504 12124
rect 14461 12087 14519 12093
rect 14461 12053 14473 12087
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 5316 11852 10425 11880
rect 5316 11840 5322 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 10413 11843 10471 11849
rect 12618 11840 12624 11892
rect 12676 11840 12682 11892
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 13906 11880 13912 11892
rect 13688 11852 13912 11880
rect 13688 11840 13694 11852
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 15562 11880 15568 11892
rect 14507 11852 15568 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 5166 11783 5172 11824
rect 5151 11777 5172 11783
rect 1486 11704 1492 11756
rect 1544 11704 1550 11756
rect 5151 11743 5163 11777
rect 5224 11772 5230 11824
rect 8846 11812 8852 11824
rect 7944 11784 8852 11812
rect 5197 11746 5212 11772
rect 6917 11747 6975 11753
rect 5197 11743 5209 11746
rect 5151 11737 5209 11743
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7374 11744 7380 11756
rect 6963 11716 7380 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 7835 11747 7893 11753
rect 7835 11713 7847 11747
rect 7881 11744 7893 11747
rect 7944 11744 7972 11784
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 9125 11815 9183 11821
rect 9125 11781 9137 11815
rect 9171 11812 9183 11815
rect 9214 11812 9220 11824
rect 9171 11784 9220 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 9493 11815 9551 11821
rect 9493 11781 9505 11815
rect 9539 11812 9551 11815
rect 10042 11812 10048 11824
rect 9539 11784 10048 11812
rect 9539 11781 9551 11784
rect 9493 11775 9551 11781
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 10226 11772 10232 11824
rect 10284 11772 10290 11824
rect 7881 11716 7972 11744
rect 9401 11747 9459 11753
rect 7881 11713 7893 11716
rect 7835 11707 7893 11713
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 9766 11744 9772 11756
rect 9447 11716 9772 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11744 9919 11747
rect 9907 11716 10640 11744
rect 9907 11713 9919 11716
rect 9861 11707 9919 11713
rect 4890 11636 4896 11688
rect 4948 11636 4954 11688
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7282 11676 7288 11688
rect 6880 11648 7288 11676
rect 6880 11636 6886 11648
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 7561 11679 7619 11685
rect 7561 11676 7573 11679
rect 7524 11648 7573 11676
rect 7524 11636 7530 11648
rect 7561 11645 7573 11648
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 8588 11648 8970 11676
rect 1026 11568 1032 11620
rect 1084 11608 1090 11620
rect 8588 11617 8616 11648
rect 8573 11611 8631 11617
rect 1084 11580 1716 11608
rect 1084 11568 1090 11580
rect 842 11500 848 11552
rect 900 11540 906 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 900 11512 1593 11540
rect 900 11500 906 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1688 11540 1716 11580
rect 5552 11580 7328 11608
rect 5552 11540 5580 11580
rect 7300 11552 7328 11580
rect 8573 11577 8585 11611
rect 8619 11577 8631 11611
rect 8573 11571 8631 11577
rect 1688 11512 5580 11540
rect 5905 11543 5963 11549
rect 1581 11503 1639 11509
rect 5905 11509 5917 11543
rect 5951 11540 5963 11543
rect 6914 11540 6920 11552
rect 5951 11512 6920 11540
rect 5951 11509 5963 11512
rect 5905 11503 5963 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 7006 11500 7012 11552
rect 7064 11500 7070 11552
rect 7282 11500 7288 11552
rect 7340 11500 7346 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 8386 11540 8392 11552
rect 7524 11512 8392 11540
rect 7524 11500 7530 11512
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 10612 11540 10640 11716
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 10744 11716 11989 11744
rect 10744 11704 10750 11716
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 12636 11744 12664 11840
rect 12636 11716 12965 11744
rect 11977 11707 12035 11713
rect 11146 11636 11152 11688
rect 11204 11636 11210 11688
rect 11698 11636 11704 11688
rect 11756 11636 11762 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 11808 11648 12633 11676
rect 11164 11608 11192 11636
rect 11808 11608 11836 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 12805 11679 12863 11685
rect 12805 11645 12817 11679
rect 12851 11645 12863 11679
rect 12937 11676 12965 11716
rect 13630 11704 13636 11756
rect 13688 11753 13694 11756
rect 13688 11747 13716 11753
rect 13704 11713 13716 11747
rect 13688 11707 13716 11713
rect 13688 11704 13694 11707
rect 13814 11704 13820 11756
rect 13872 11704 13878 11756
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 12937 11648 13553 11676
rect 12805 11639 12863 11645
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 12820 11608 12848 11639
rect 11164 11580 11836 11608
rect 12268 11580 12848 11608
rect 12268 11552 12296 11580
rect 13262 11568 13268 11620
rect 13320 11568 13326 11620
rect 12250 11540 12256 11552
rect 10612 11512 12256 11540
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 7466 11336 7472 11348
rect 6472 11308 7472 11336
rect 4890 11160 4896 11212
rect 4948 11200 4954 11212
rect 5261 11203 5319 11209
rect 5261 11200 5273 11203
rect 4948 11172 5273 11200
rect 4948 11160 4954 11172
rect 5261 11169 5273 11172
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 5535 11135 5593 11141
rect 5535 11101 5547 11135
rect 5581 11132 5593 11135
rect 6472 11132 6500 11308
rect 7466 11296 7472 11308
rect 7524 11296 7530 11348
rect 8754 11336 8760 11348
rect 7576 11308 8760 11336
rect 7576 11268 7604 11308
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9858 11336 9864 11348
rect 8904 11308 9864 11336
rect 8904 11296 8910 11308
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 10042 11296 10048 11348
rect 10100 11296 10106 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 13081 11339 13139 11345
rect 10928 11308 13032 11336
rect 10928 11296 10934 11308
rect 7116 11240 7604 11268
rect 8864 11268 8892 11296
rect 9876 11268 9904 11296
rect 11146 11268 11152 11280
rect 8864 11240 9076 11268
rect 9876 11240 11152 11268
rect 6822 11200 6828 11212
rect 6806 11160 6828 11200
rect 6880 11160 6886 11212
rect 5581 11104 6500 11132
rect 5581 11101 5593 11104
rect 5535 11095 5593 11101
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 6806 11132 6834 11160
rect 7116 11141 7144 11240
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 9048 11209 9076 11240
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 11238 11228 11244 11280
rect 11296 11228 11302 11280
rect 13004 11268 13032 11308
rect 13081 11305 13093 11339
rect 13127 11336 13139 11339
rect 13262 11336 13268 11348
rect 13127 11308 13268 11336
rect 13127 11305 13139 11308
rect 13081 11299 13139 11305
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13906 11296 13912 11348
rect 13964 11296 13970 11348
rect 14458 11296 14464 11348
rect 14516 11296 14522 11348
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 13004 11240 13645 11268
rect 13633 11237 13645 11240
rect 13679 11237 13691 11271
rect 13633 11231 13691 11237
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7524 11172 7573 11200
rect 7524 11160 7530 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 7561 11163 7619 11169
rect 7975 11203 8033 11209
rect 7975 11169 7987 11203
rect 8021 11200 8033 11203
rect 9033 11203 9091 11209
rect 8021 11172 8984 11200
rect 8021 11169 8033 11172
rect 7975 11163 8033 11169
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6604 11104 6929 11132
rect 6604 11092 6610 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 7834 11092 7840 11144
rect 7892 11092 7898 11144
rect 8110 11092 8116 11144
rect 8168 11092 8174 11144
rect 8956 11076 8984 11172
rect 9033 11169 9045 11203
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 10226 11160 10232 11212
rect 10284 11160 10290 11212
rect 11256 11200 11284 11228
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 11256 11172 11437 11200
rect 11425 11169 11437 11172
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 11882 11160 11888 11212
rect 11940 11160 11946 11212
rect 14642 11200 14648 11212
rect 13464 11172 14648 11200
rect 9306 11092 9312 11144
rect 9364 11092 9370 11144
rect 1489 11067 1547 11073
rect 1489 11033 1501 11067
rect 1535 11064 1547 11067
rect 2406 11064 2412 11076
rect 1535 11036 2412 11064
rect 1535 11033 1547 11036
rect 1489 11027 1547 11033
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 3878 11024 3884 11076
rect 3936 11064 3942 11076
rect 4982 11064 4988 11076
rect 3936 11036 4988 11064
rect 3936 11024 3942 11036
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 8588 11036 8892 11064
rect 1578 10956 1584 11008
rect 1636 10956 1642 11008
rect 6273 10999 6331 11005
rect 6273 10965 6285 10999
rect 6319 10996 6331 10999
rect 6454 10996 6460 11008
rect 6319 10968 6460 10996
rect 6319 10965 6331 10968
rect 6273 10959 6331 10965
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 6638 10956 6644 11008
rect 6696 10956 6702 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 8588 10996 8616 11036
rect 6788 10968 8616 10996
rect 6788 10956 6794 10968
rect 8754 10956 8760 11008
rect 8812 10956 8818 11008
rect 8864 10996 8892 11036
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 10244 11064 10272 11160
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11054 11132 11060 11144
rect 10919 11104 11060 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11132 11207 11135
rect 11900 11132 11928 11160
rect 11195 11104 11928 11132
rect 11195 11101 11207 11104
rect 11149 11095 11207 11101
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 13464 11141 13492 11172
rect 14642 11160 14648 11172
rect 14700 11160 14706 11212
rect 12069 11135 12127 11141
rect 12069 11132 12081 11135
rect 12032 11104 12081 11132
rect 12032 11092 12038 11104
rect 12069 11101 12081 11104
rect 12115 11101 12127 11135
rect 12311 11135 12369 11141
rect 12311 11132 12323 11135
rect 12069 11095 12127 11101
rect 12176 11104 12323 11132
rect 11606 11064 11612 11076
rect 8996 11036 10272 11064
rect 11072 11036 11612 11064
rect 8996 11024 9002 11036
rect 10594 10996 10600 11008
rect 8864 10968 10600 10996
rect 10594 10956 10600 10968
rect 10652 10956 10658 11008
rect 11072 11005 11100 11036
rect 11606 11024 11612 11036
rect 11664 11024 11670 11076
rect 11057 10999 11115 11005
rect 11057 10965 11069 10999
rect 11103 10965 11115 10999
rect 12084 10996 12112 11095
rect 12176 11076 12204 11104
rect 12311 11101 12323 11104
rect 12357 11101 12369 11135
rect 12311 11095 12369 11101
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14182 11132 14188 11144
rect 13771 11104 14188 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 15102 11132 15108 11144
rect 14323 11104 15108 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 12158 11024 12164 11076
rect 12216 11024 12222 11076
rect 12710 10996 12716 11008
rect 12084 10968 12716 10996
rect 11057 10959 11115 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 15838 10888 15844 10940
rect 15896 10888 15902 10940
rect 1104 10832 14971 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1544 10764 1593 10792
rect 1544 10752 1550 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 7006 10792 7012 10804
rect 1581 10755 1639 10761
rect 5828 10764 7012 10792
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 1811 10628 2774 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 2746 10452 2774 10628
rect 5828 10588 5856 10764
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 7742 10792 7748 10804
rect 7616 10764 7748 10792
rect 7616 10752 7622 10764
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 10836 10764 11910 10792
rect 10836 10752 10842 10764
rect 6730 10724 6736 10736
rect 6564 10696 6736 10724
rect 6564 10665 6592 10696
rect 6730 10684 6736 10696
rect 6788 10684 6794 10736
rect 11790 10684 11796 10736
rect 11848 10684 11854 10736
rect 11882 10724 11910 10764
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12158 10792 12164 10804
rect 12032 10764 12164 10792
rect 12032 10752 12038 10764
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 13814 10752 13820 10804
rect 13872 10752 13878 10804
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 15856 10792 15884 10888
rect 14415 10764 15884 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 14384 10724 14412 10755
rect 11882 10696 14412 10724
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 6549 10659 6607 10665
rect 5951 10628 6500 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 6472 10600 6500 10628
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 6696 10628 6960 10656
rect 6696 10616 6702 10628
rect 5997 10591 6055 10597
rect 5997 10588 6009 10591
rect 5828 10560 6009 10588
rect 5997 10557 6009 10560
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10557 6239 10591
rect 6181 10551 6239 10557
rect 6196 10520 6224 10551
rect 6454 10548 6460 10600
rect 6512 10548 6518 10600
rect 6733 10591 6791 10597
rect 6733 10557 6745 10591
rect 6779 10588 6791 10591
rect 6822 10588 6828 10600
rect 6779 10560 6828 10588
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 6932 10588 6960 10628
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 8478 10616 8484 10668
rect 8536 10656 8542 10668
rect 9306 10656 9312 10668
rect 8536 10628 9312 10656
rect 8536 10616 8542 10628
rect 9306 10616 9312 10628
rect 9364 10656 9370 10668
rect 11808 10656 11836 10684
rect 9364 10628 11836 10656
rect 9364 10616 9370 10628
rect 11808 10597 11836 10628
rect 12342 10616 12348 10668
rect 12400 10656 12406 10668
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 12400 10628 12449 10656
rect 12400 10616 12406 10628
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 13047 10659 13105 10665
rect 13047 10656 13059 10659
rect 12437 10619 12495 10625
rect 12636 10628 13059 10656
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 6932 10560 7481 10588
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7607 10591 7665 10597
rect 7607 10557 7619 10591
rect 7653 10588 7665 10591
rect 8665 10591 8723 10597
rect 8665 10588 8677 10591
rect 7653 10560 8677 10588
rect 7653 10557 7665 10560
rect 7607 10551 7665 10557
rect 8665 10557 8677 10560
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 6196 10492 6868 10520
rect 6840 10464 6868 10492
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7193 10523 7251 10529
rect 7193 10520 7205 10523
rect 6972 10492 7205 10520
rect 6972 10480 6978 10492
rect 7193 10489 7205 10492
rect 7239 10489 7251 10523
rect 7193 10483 7251 10489
rect 4154 10452 4160 10464
rect 2746 10424 4160 10452
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 6089 10455 6147 10461
rect 6089 10452 6101 10455
rect 4304 10424 6101 10452
rect 4304 10412 4310 10424
rect 6089 10421 6101 10424
rect 6135 10421 6147 10455
rect 6089 10415 6147 10421
rect 6822 10412 6828 10464
rect 6880 10412 6886 10464
rect 7208 10452 7236 10483
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 11238 10520 11244 10532
rect 10744 10492 11244 10520
rect 10744 10480 10750 10492
rect 11238 10480 11244 10492
rect 11296 10480 11302 10532
rect 11532 10520 11560 10551
rect 12158 10548 12164 10600
rect 12216 10588 12222 10600
rect 12636 10588 12664 10628
rect 13047 10625 13059 10628
rect 13093 10625 13105 10659
rect 13047 10619 13105 10625
rect 14182 10616 14188 10668
rect 14240 10616 14246 10668
rect 12216 10560 12664 10588
rect 12216 10548 12222 10560
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12768 10560 12817 10588
rect 12768 10548 12774 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 11532 10492 12940 10520
rect 7466 10452 7472 10464
rect 7208 10424 7472 10452
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 12434 10452 12440 10464
rect 11756 10424 12440 10452
rect 11756 10412 11762 10424
rect 12434 10412 12440 10424
rect 12492 10452 12498 10464
rect 12621 10455 12679 10461
rect 12621 10452 12633 10455
rect 12492 10424 12633 10452
rect 12492 10412 12498 10424
rect 12621 10421 12633 10424
rect 12667 10421 12679 10455
rect 12912 10452 12940 10492
rect 15470 10452 15476 10464
rect 12912 10424 15476 10452
rect 12621 10415 12679 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 2406 10208 2412 10260
rect 2464 10208 2470 10260
rect 6822 10208 6828 10260
rect 6880 10208 6886 10260
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7432 10220 7849 10248
rect 7432 10208 7438 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 8386 10208 8392 10260
rect 8444 10208 8450 10260
rect 10318 10208 10324 10260
rect 10376 10208 10382 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11112 10220 11989 10248
rect 11112 10208 11118 10220
rect 11977 10217 11989 10220
rect 12023 10248 12035 10251
rect 12250 10248 12256 10260
rect 12023 10220 12256 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12250 10208 12256 10220
rect 12308 10248 12314 10260
rect 12618 10248 12624 10260
rect 12308 10220 12624 10248
rect 12308 10208 12314 10220
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 12986 10248 12992 10260
rect 12768 10220 12992 10248
rect 12768 10208 12774 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13630 10208 13636 10260
rect 13688 10208 13694 10260
rect 13909 10251 13967 10257
rect 13909 10217 13921 10251
rect 13955 10248 13967 10251
rect 13998 10248 14004 10260
rect 13955 10220 14004 10248
rect 13955 10217 13967 10220
rect 13909 10211 13967 10217
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 2225 10183 2283 10189
rect 2225 10149 2237 10183
rect 2271 10180 2283 10183
rect 3970 10180 3976 10192
rect 2271 10152 3976 10180
rect 2271 10149 2283 10152
rect 2225 10143 2283 10149
rect 3970 10140 3976 10152
rect 4028 10140 4034 10192
rect 7561 10183 7619 10189
rect 7561 10149 7573 10183
rect 7607 10149 7619 10183
rect 7561 10143 7619 10149
rect 1026 10004 1032 10056
rect 1084 10044 1090 10056
rect 2041 10047 2099 10053
rect 2041 10044 2053 10047
rect 1084 10016 2053 10044
rect 1084 10004 1090 10016
rect 2041 10013 2053 10016
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2363 10016 6408 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 1489 9979 1547 9985
rect 1489 9945 1501 9979
rect 1535 9976 1547 9979
rect 2774 9976 2780 9988
rect 1535 9948 2780 9976
rect 1535 9945 1547 9948
rect 1489 9939 1547 9945
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 6380 9976 6408 10016
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 6512 10016 6745 10044
rect 6512 10004 6518 10016
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 7576 10044 7604 10143
rect 8404 10112 8432 10208
rect 10336 10180 10364 10208
rect 10060 10152 10364 10180
rect 13648 10180 13676 10208
rect 14461 10183 14519 10189
rect 14461 10180 14473 10183
rect 13648 10152 14473 10180
rect 7760 10084 8432 10112
rect 7760 10053 7788 10084
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 10060 10121 10088 10152
rect 14461 10149 14473 10152
rect 14507 10149 14519 10183
rect 14461 10143 14519 10149
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9732 10084 10057 10112
rect 9732 10072 9738 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10284 10084 10517 10112
rect 10284 10072 10290 10084
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10594 10072 10600 10124
rect 10652 10112 10658 10124
rect 10898 10115 10956 10121
rect 10898 10112 10910 10115
rect 10652 10084 10910 10112
rect 10652 10072 10658 10084
rect 10898 10081 10910 10084
rect 10944 10081 10956 10115
rect 10898 10075 10956 10081
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 11238 10112 11244 10124
rect 11103 10084 11244 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 11664 10084 12081 10112
rect 11664 10072 11670 10084
rect 12069 10081 12081 10084
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 12710 10072 12716 10124
rect 12768 10072 12774 10124
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12860 10084 13001 10112
rect 12860 10072 12866 10084
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13127 10115 13185 10121
rect 13127 10081 13139 10115
rect 13173 10112 13185 10115
rect 13446 10112 13452 10124
rect 13173 10084 13452 10112
rect 13173 10081 13185 10084
rect 13127 10075 13185 10081
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 6963 10016 7604 10044
rect 7745 10047 7803 10053
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8754 10044 8760 10056
rect 8067 10016 8760 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 9861 10047 9919 10053
rect 9861 10044 9873 10047
rect 9646 10016 9873 10044
rect 6638 9976 6644 9988
rect 6380 9948 6644 9976
rect 6638 9936 6644 9948
rect 6696 9936 6702 9988
rect 9306 9936 9312 9988
rect 9364 9976 9370 9988
rect 9490 9976 9496 9988
rect 9364 9948 9496 9976
rect 9364 9936 9370 9948
rect 9490 9936 9496 9948
rect 9548 9976 9554 9988
rect 9646 9976 9674 10016
rect 9861 10013 9873 10016
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 10778 10004 10784 10056
rect 10836 10004 10842 10056
rect 11790 10004 11796 10056
rect 11848 10004 11854 10056
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12268 9976 12296 10007
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 9548 9948 9674 9976
rect 11624 9948 12296 9976
rect 9548 9936 9554 9948
rect 11624 9920 11652 9948
rect 14274 9936 14280 9988
rect 14332 9936 14338 9988
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 10962 9908 10968 9920
rect 4212 9880 10968 9908
rect 4212 9868 4218 9880
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11606 9868 11612 9920
rect 11664 9868 11670 9920
rect 11701 9911 11759 9917
rect 11701 9877 11713 9911
rect 11747 9908 11759 9911
rect 11974 9908 11980 9920
rect 11747 9880 11980 9908
rect 11747 9877 11759 9880
rect 11701 9871 11759 9877
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 12710 9908 12716 9920
rect 12308 9880 12716 9908
rect 12308 9868 12314 9880
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 2774 9664 2780 9716
rect 2832 9664 2838 9716
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10778 9704 10784 9716
rect 10468 9676 10784 9704
rect 10468 9664 10474 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 13446 9704 13452 9716
rect 11020 9676 13452 9704
rect 11020 9664 11026 9676
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6604 9608 7144 9636
rect 6604 9596 6610 9608
rect 7116 9580 7144 9608
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 7650 9636 7656 9648
rect 7432 9608 7656 9636
rect 7432 9596 7438 9608
rect 7650 9596 7656 9608
rect 7708 9636 7714 9648
rect 7708 9608 9720 9636
rect 7708 9596 7714 9608
rect 9692 9580 9720 9608
rect 11606 9596 11612 9648
rect 11664 9596 11670 9648
rect 1671 9571 1729 9577
rect 1671 9537 1683 9571
rect 1717 9568 1729 9571
rect 1762 9568 1768 9580
rect 1717 9540 1768 9568
rect 1717 9537 1729 9540
rect 1671 9531 1729 9537
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2424 9540 2973 9568
rect 1394 9460 1400 9512
rect 1452 9460 1458 9512
rect 2424 9441 2452 9540
rect 2961 9537 2973 9540
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 6454 9528 6460 9580
rect 6512 9528 6518 9580
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6914 9568 6920 9580
rect 6687 9540 6920 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7098 9528 7104 9580
rect 7156 9528 7162 9580
rect 9490 9528 9496 9580
rect 9548 9528 9554 9580
rect 9674 9528 9680 9580
rect 9732 9528 9738 9580
rect 10410 9528 10416 9580
rect 10468 9528 10474 9580
rect 10594 9577 10600 9580
rect 10551 9571 10600 9577
rect 10551 9537 10563 9571
rect 10597 9537 10600 9571
rect 10551 9531 10600 9537
rect 10594 9528 10600 9531
rect 10652 9528 10658 9580
rect 11624 9568 11652 9596
rect 11440 9566 11652 9568
rect 11701 9571 11759 9577
rect 11701 9566 11713 9571
rect 11440 9540 11713 9566
rect 11440 9512 11468 9540
rect 11624 9538 11713 9540
rect 11701 9537 11713 9538
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 12526 9528 12532 9580
rect 12584 9577 12590 9580
rect 12584 9571 12633 9577
rect 12584 9537 12587 9571
rect 12621 9537 12633 9571
rect 12584 9531 12633 9537
rect 12584 9528 12590 9531
rect 12710 9528 12716 9580
rect 12768 9528 12774 9580
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 13280 9540 13921 9568
rect 8294 9460 8300 9512
rect 8352 9500 8358 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 8352 9472 8401 9500
rect 8352 9460 8358 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 10042 9500 10048 9512
rect 8389 9463 8447 9469
rect 9968 9472 10048 9500
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9401 2467 9435
rect 2409 9395 2467 9401
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 8938 9432 8944 9444
rect 7524 9404 8944 9432
rect 7524 9392 7530 9404
rect 8938 9392 8944 9404
rect 8996 9432 9002 9444
rect 9858 9432 9864 9444
rect 8996 9404 9864 9432
rect 8996 9392 9002 9404
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 9968 9364 9996 9472
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9500 10747 9503
rect 10870 9500 10876 9512
rect 10735 9472 10876 9500
rect 10735 9469 10747 9472
rect 10689 9463 10747 9469
rect 10870 9460 10876 9472
rect 10928 9500 10934 9512
rect 11238 9500 11244 9512
rect 10928 9472 11244 9500
rect 10928 9460 10934 9472
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 11422 9460 11428 9512
rect 11480 9460 11486 9512
rect 11514 9460 11520 9512
rect 11572 9460 11578 9512
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 13280 9500 13308 9540
rect 13909 9537 13921 9540
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 12492 9472 13308 9500
rect 13633 9503 13691 9509
rect 12492 9460 12498 9472
rect 13633 9469 13645 9503
rect 13679 9500 13691 9503
rect 13814 9500 13820 9512
rect 13679 9472 13820 9500
rect 13679 9469 13691 9472
rect 13633 9463 13691 9469
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 10137 9435 10195 9441
rect 10137 9401 10149 9435
rect 10183 9401 10195 9435
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 10137 9395 10195 9401
rect 11072 9404 12173 9432
rect 7892 9336 9996 9364
rect 7892 9324 7898 9336
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10152 9364 10180 9395
rect 11072 9364 11100 9404
rect 12161 9401 12173 9404
rect 12207 9401 12219 9435
rect 12161 9395 12219 9401
rect 10100 9336 11100 9364
rect 10100 9324 10106 9336
rect 11330 9324 11336 9376
rect 11388 9324 11394 9376
rect 13354 9324 13360 9376
rect 13412 9324 13418 9376
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 1118 9120 1124 9172
rect 1176 9160 1182 9172
rect 1176 9132 2774 9160
rect 1176 9120 1182 9132
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 2746 8956 2774 9132
rect 6454 9120 6460 9172
rect 6512 9120 6518 9172
rect 6546 9120 6552 9172
rect 6604 9120 6610 9172
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6696 9132 6745 9160
rect 6696 9120 6702 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 8018 9120 8024 9172
rect 8076 9160 8082 9172
rect 8076 9132 9628 9160
rect 8076 9120 8082 9132
rect 6181 9095 6239 9101
rect 6181 9061 6193 9095
rect 6227 9092 6239 9095
rect 6472 9092 6500 9120
rect 6227 9064 6500 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 4890 8984 4896 9036
rect 4948 9024 4954 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 4948 8996 5181 9024
rect 4948 8984 4954 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 6472 8956 6500 9064
rect 6564 9024 6592 9120
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 8938 9092 8944 9104
rect 8628 9064 8944 9092
rect 8628 9052 8634 9064
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 6825 9027 6883 9033
rect 6825 9024 6837 9027
rect 6564 8996 6837 9024
rect 6825 8993 6837 8996
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7466 9024 7472 9036
rect 6963 8996 7472 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 9024 7619 9027
rect 7650 9024 7656 9036
rect 7607 8996 7656 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 8018 9033 8024 9036
rect 7975 9027 8024 9033
rect 7975 8993 7987 9027
rect 8021 8993 8024 9027
rect 7975 8987 8024 8993
rect 8018 8984 8024 8987
rect 8076 8984 8082 9036
rect 8113 9027 8171 9033
rect 8113 8993 8125 9027
rect 8159 9024 8171 9027
rect 8478 9024 8484 9036
rect 8159 8996 8484 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 9600 8968 9628 9132
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10502 9160 10508 9172
rect 10192 9132 10508 9160
rect 10192 9120 10198 9132
rect 10502 9120 10508 9132
rect 10560 9160 10566 9172
rect 11054 9160 11060 9172
rect 10560 9132 11060 9160
rect 10560 9120 10566 9132
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11330 9120 11336 9172
rect 11388 9120 11394 9172
rect 13354 9120 13360 9172
rect 13412 9120 13418 9172
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 13504 9132 14381 9160
rect 13504 9120 13510 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 14369 9123 14427 9129
rect 9858 8984 9864 9036
rect 9916 8984 9922 9036
rect 10318 9033 10324 9036
rect 10275 9027 10324 9033
rect 10275 8993 10287 9027
rect 10321 8993 10324 9027
rect 10275 8987 10324 8993
rect 10318 8984 10324 8987
rect 10376 8984 10382 9036
rect 10413 9027 10471 9033
rect 10413 8993 10425 9027
rect 10459 9024 10471 9027
rect 10962 9024 10968 9036
rect 10459 8996 10968 9024
rect 10459 8993 10471 8996
rect 10413 8987 10471 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11348 9024 11376 9120
rect 11790 9052 11796 9104
rect 11848 9052 11854 9104
rect 12069 9027 12127 9033
rect 12069 9024 12081 9027
rect 11348 8996 12081 9024
rect 12069 8993 12081 8996
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 12207 9027 12265 9033
rect 12207 8993 12219 9027
rect 12253 9024 12265 9027
rect 13372 9024 13400 9120
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 13909 9095 13967 9101
rect 13909 9092 13921 9095
rect 13596 9064 13921 9092
rect 13596 9052 13602 9064
rect 13909 9061 13921 9064
rect 13955 9061 13967 9095
rect 13909 9055 13967 9061
rect 12253 8996 13400 9024
rect 12253 8993 12265 8996
rect 12207 8987 12265 8993
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 1655 8929 1713 8935
rect 1655 8895 1667 8929
rect 1701 8926 1713 8929
rect 2746 8929 5488 8956
rect 2746 8928 5439 8929
rect 1701 8895 1716 8926
rect 1655 8889 1716 8895
rect 1688 8888 1716 8889
rect 1854 8888 1860 8900
rect 1688 8860 1860 8888
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 5427 8895 5439 8928
rect 5473 8895 5488 8929
rect 6472 8928 6561 8956
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 7098 8916 7104 8968
rect 7156 8916 7162 8968
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8812 8928 9137 8956
rect 8812 8916 8818 8928
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9398 8916 9404 8968
rect 9456 8916 9462 8968
rect 9582 8916 9588 8968
rect 9640 8916 9646 8968
rect 10134 8916 10140 8968
rect 10192 8965 10198 8968
rect 10192 8959 10213 8965
rect 10201 8925 10213 8959
rect 10192 8919 10213 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 11149 8959 11207 8965
rect 11149 8956 11161 8959
rect 11103 8928 11161 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 11149 8925 11161 8928
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 10192 8916 10198 8919
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 11296 8928 11345 8956
rect 11296 8916 11302 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 12342 8916 12348 8968
rect 12400 8916 12406 8968
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13648 8956 13676 8984
rect 13035 8928 13676 8956
rect 14277 8959 14335 8965
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 15102 8956 15108 8968
rect 14323 8928 15108 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 5427 8889 5488 8895
rect 5460 8832 5488 8889
rect 13354 8848 13360 8900
rect 13412 8848 13418 8900
rect 13722 8848 13728 8900
rect 13780 8848 13786 8900
rect 2406 8780 2412 8832
rect 2464 8780 2470 8832
rect 5442 8780 5448 8832
rect 5500 8780 5506 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 8757 8823 8815 8829
rect 8757 8820 8769 8823
rect 7524 8792 8769 8820
rect 7524 8780 7530 8792
rect 8757 8789 8769 8792
rect 8803 8789 8815 8823
rect 8757 8783 8815 8789
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 10042 8820 10048 8832
rect 9916 8792 10048 8820
rect 9916 8780 9922 8792
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 13446 8820 13452 8832
rect 11756 8792 13452 8820
rect 11756 8780 11762 8792
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1504 8588 1961 8616
rect 1504 8557 1532 8588
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 1949 8579 2007 8585
rect 2406 8576 2412 8628
rect 2464 8576 2470 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 6549 8619 6607 8625
rect 6549 8585 6561 8619
rect 6595 8616 6607 8619
rect 6638 8616 6644 8628
rect 6595 8588 6644 8616
rect 6595 8585 6607 8588
rect 6549 8579 6607 8585
rect 1489 8551 1547 8557
rect 1489 8517 1501 8551
rect 1535 8517 1547 8551
rect 1489 8511 1547 8517
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2424 8480 2452 8576
rect 6012 8548 6040 8579
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 6914 8576 6920 8628
rect 6972 8576 6978 8628
rect 7466 8576 7472 8628
rect 7524 8576 7530 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 7576 8588 9229 8616
rect 7484 8548 7512 8576
rect 6012 8520 6500 8548
rect 6472 8489 6500 8520
rect 7024 8520 7512 8548
rect 2179 8452 2452 8480
rect 6181 8483 6239 8489
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6457 8483 6515 8489
rect 6457 8449 6469 8483
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 6196 8412 6224 8443
rect 7024 8412 7052 8520
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 7576 8480 7604 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9582 8616 9588 8628
rect 9217 8579 9275 8585
rect 9508 8588 9588 8616
rect 7147 8452 7604 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 8294 8440 8300 8492
rect 8352 8440 8358 8492
rect 9508 8489 9536 8588
rect 9582 8576 9588 8588
rect 9640 8616 9646 8628
rect 11606 8616 11612 8628
rect 9640 8588 11612 8616
rect 9640 8576 9646 8588
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 11790 8576 11796 8628
rect 11848 8616 11854 8628
rect 12529 8619 12587 8625
rect 12529 8616 12541 8619
rect 11848 8588 12541 8616
rect 11848 8576 11854 8588
rect 12529 8585 12541 8588
rect 12575 8585 12587 8619
rect 12986 8616 12992 8628
rect 12529 8579 12587 8585
rect 12728 8588 12992 8616
rect 12434 8548 12440 8560
rect 11440 8520 12440 8548
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 9723 8452 9812 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 9784 8424 9812 8452
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10502 8440 10508 8492
rect 10560 8489 10566 8492
rect 10560 8483 10588 8489
rect 10576 8449 10588 8483
rect 10560 8443 10588 8449
rect 10560 8440 10566 8443
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 6196 8384 7052 8412
rect 7190 8372 7196 8424
rect 7248 8372 7254 8424
rect 7374 8372 7380 8424
rect 7432 8372 7438 8424
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8381 7619 8415
rect 8435 8415 8493 8421
rect 8435 8412 8447 8415
rect 7561 8375 7619 8381
rect 8128 8384 8447 8412
rect 1670 8304 1676 8356
rect 1728 8304 1734 8356
rect 7208 8344 7236 8372
rect 7576 8344 7604 8375
rect 7208 8316 7604 8344
rect 7650 8304 7656 8356
rect 7708 8344 7714 8356
rect 8021 8347 8079 8353
rect 8021 8344 8033 8347
rect 7708 8316 8033 8344
rect 7708 8304 7714 8316
rect 8021 8313 8033 8316
rect 8067 8313 8079 8347
rect 8021 8307 8079 8313
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 8128 8276 8156 8384
rect 8435 8381 8447 8384
rect 8481 8381 8493 8415
rect 8435 8375 8493 8381
rect 8583 8415 8641 8421
rect 8583 8381 8595 8415
rect 8629 8412 8641 8415
rect 8629 8384 8984 8412
rect 8629 8381 8641 8384
rect 8583 8375 8641 8381
rect 7984 8248 8156 8276
rect 7984 8236 7990 8248
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 8956 8276 8984 8384
rect 9766 8372 9772 8424
rect 9824 8372 9830 8424
rect 9876 8412 9904 8440
rect 10413 8415 10471 8421
rect 10413 8412 10425 8415
rect 9876 8384 10425 8412
rect 10413 8381 10425 8384
rect 10459 8412 10471 8415
rect 11440 8412 11468 8520
rect 12434 8508 12440 8520
rect 12492 8508 12498 8560
rect 11791 8483 11849 8489
rect 11791 8449 11803 8483
rect 11837 8480 11849 8483
rect 11882 8480 11888 8492
rect 11837 8452 11888 8480
rect 11837 8449 11849 8452
rect 11791 8443 11849 8449
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 10459 8384 11468 8412
rect 11517 8415 11575 8421
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 11517 8381 11529 8415
rect 11563 8381 11575 8415
rect 12728 8412 12756 8588
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13906 8576 13912 8628
rect 13964 8576 13970 8628
rect 12802 8508 12808 8560
rect 12860 8548 12866 8560
rect 12860 8520 13124 8548
rect 12860 8508 12866 8520
rect 13096 8510 13124 8520
rect 13155 8513 13213 8519
rect 13155 8510 13167 8513
rect 13096 8482 13167 8510
rect 13155 8479 13167 8482
rect 13201 8479 13213 8513
rect 13155 8473 13213 8479
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 11517 8375 11575 8381
rect 12544 8384 12909 8412
rect 9784 8344 9812 8372
rect 8536 8248 8984 8276
rect 9692 8316 9812 8344
rect 9692 8276 9720 8316
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 10137 8347 10195 8353
rect 10137 8344 10149 8347
rect 9916 8316 10149 8344
rect 9916 8304 9922 8316
rect 10137 8313 10149 8316
rect 10183 8344 10195 8347
rect 10226 8344 10232 8356
rect 10183 8316 10232 8344
rect 10183 8313 10195 8316
rect 10137 8307 10195 8313
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 11330 8304 11336 8356
rect 11388 8304 11394 8356
rect 11422 8304 11428 8356
rect 11480 8344 11486 8356
rect 11532 8344 11560 8375
rect 11480 8316 11560 8344
rect 11480 8304 11486 8316
rect 10870 8276 10876 8288
rect 9692 8248 10876 8276
rect 8536 8236 8542 8248
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 12544 8276 12572 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 11112 8248 12572 8276
rect 11112 8236 11118 8248
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 12894 8276 12900 8288
rect 12676 8248 12900 8276
rect 12676 8236 12682 8248
rect 12894 8236 12900 8248
rect 12952 8276 12958 8288
rect 13814 8276 13820 8288
rect 12952 8248 13820 8276
rect 12952 8236 12958 8248
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7708 8044 7849 8072
rect 7708 8032 7714 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 7926 8032 7932 8084
rect 7984 8072 7990 8084
rect 8754 8072 8760 8084
rect 7984 8044 8760 8072
rect 7984 8032 7990 8044
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 11940 8044 12296 8072
rect 11940 8032 11946 8044
rect 12268 8004 12296 8044
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12400 8044 12633 8072
rect 12400 8032 12406 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 13814 8032 13820 8084
rect 13872 8032 13878 8084
rect 13906 8004 13912 8016
rect 12268 7976 13912 8004
rect 13906 7964 13912 7976
rect 13964 8004 13970 8016
rect 14461 8007 14519 8013
rect 14461 8004 14473 8007
rect 13964 7976 14473 8004
rect 13964 7964 13970 7976
rect 14461 7973 14473 7976
rect 14507 7973 14519 8007
rect 14461 7967 14519 7973
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 4948 7908 6837 7936
rect 4948 7896 4954 7908
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7936 10747 7939
rect 11514 7936 11520 7948
rect 10735 7908 11520 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 1486 7760 1492 7812
rect 1544 7760 1550 7812
rect 6840 7800 6868 7899
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 7083 7841 7141 7847
rect 6914 7800 6920 7812
rect 6840 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 7083 7807 7095 7841
rect 7129 7838 7141 7841
rect 7129 7807 7144 7838
rect 10870 7828 10876 7880
rect 10928 7868 10934 7880
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10928 7840 10977 7868
rect 10928 7828 10934 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 11606 7868 11612 7880
rect 11480 7840 11612 7868
rect 11480 7828 11486 7840
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 11883 7871 11941 7877
rect 11883 7837 11895 7871
rect 11929 7868 11941 7871
rect 12250 7868 12256 7880
rect 11929 7840 12256 7868
rect 11929 7837 11941 7840
rect 11883 7831 11941 7837
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 7083 7801 7144 7807
rect 7116 7800 7144 7801
rect 8386 7800 8392 7812
rect 7116 7772 8392 7800
rect 8386 7760 8392 7772
rect 8444 7800 8450 7812
rect 12618 7800 12624 7812
rect 8444 7772 12624 7800
rect 8444 7760 8450 7772
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 13725 7803 13783 7809
rect 13725 7769 13737 7803
rect 13771 7800 13783 7803
rect 15102 7800 15108 7812
rect 13771 7772 15108 7800
rect 13771 7769 13783 7772
rect 13725 7763 13783 7769
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 900 7704 1593 7732
rect 900 7692 906 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 1581 7695 1639 7701
rect 9398 7692 9404 7744
rect 9456 7732 9462 7744
rect 13630 7732 13636 7744
rect 9456 7704 13636 7732
rect 9456 7692 9462 7704
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 6546 7528 6552 7540
rect 5684 7500 6552 7528
rect 5684 7488 5690 7500
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 8757 7531 8815 7537
rect 8757 7497 8769 7531
rect 8803 7528 8815 7531
rect 10686 7528 10692 7540
rect 8803 7500 10692 7528
rect 8803 7497 8815 7500
rect 8757 7491 8815 7497
rect 10686 7488 10692 7500
rect 10744 7528 10750 7540
rect 10962 7528 10968 7540
rect 10744 7500 10968 7528
rect 10744 7488 10750 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11146 7488 11152 7540
rect 11204 7528 11210 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 11204 7500 11345 7528
rect 11204 7488 11210 7500
rect 11333 7497 11345 7500
rect 11379 7497 11391 7531
rect 11333 7491 11391 7497
rect 12529 7531 12587 7537
rect 12529 7497 12541 7531
rect 12575 7528 12587 7531
rect 13170 7528 13176 7540
rect 12575 7500 13176 7528
rect 12575 7497 12587 7500
rect 12529 7491 12587 7497
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 13630 7528 13636 7540
rect 13280 7500 13636 7528
rect 13081 7463 13139 7469
rect 13081 7429 13093 7463
rect 13127 7460 13139 7463
rect 13280 7460 13308 7500
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 14366 7488 14372 7540
rect 14424 7488 14430 7540
rect 13127 7432 13308 7460
rect 13357 7463 13415 7469
rect 13127 7429 13139 7432
rect 13081 7423 13139 7429
rect 13357 7429 13369 7463
rect 13403 7460 13415 7463
rect 13538 7460 13544 7472
rect 13403 7432 13544 7460
rect 13403 7429 13415 7432
rect 13357 7423 13415 7429
rect 13538 7420 13544 7432
rect 13596 7420 13602 7472
rect 13998 7460 14004 7472
rect 13832 7432 14004 7460
rect 1671 7395 1729 7401
rect 1671 7361 1683 7395
rect 1717 7392 1729 7395
rect 7006 7392 7012 7404
rect 1717 7364 7012 7392
rect 1717 7361 1729 7364
rect 1671 7355 1729 7361
rect 7006 7352 7012 7364
rect 7064 7392 7070 7404
rect 7987 7395 8045 7401
rect 7987 7392 7999 7395
rect 7064 7364 7999 7392
rect 7064 7352 7070 7364
rect 7987 7361 7999 7364
rect 8033 7361 8045 7395
rect 7987 7355 8045 7361
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 9088 7364 9505 7392
rect 9088 7352 9094 7364
rect 9493 7361 9505 7364
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 10686 7352 10692 7404
rect 10744 7352 10750 7404
rect 11790 7392 11796 7404
rect 11751 7364 11796 7392
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 13446 7352 13452 7404
rect 13504 7352 13510 7404
rect 13832 7401 13860 7432
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 14185 7463 14243 7469
rect 14185 7429 14197 7463
rect 14231 7429 14243 7463
rect 14185 7423 14243 7429
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14200 7392 14228 7423
rect 13964 7364 14228 7392
rect 13964 7352 13970 7364
rect 1394 7284 1400 7336
rect 1452 7284 1458 7336
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7650 7324 7656 7336
rect 6972 7296 7656 7324
rect 6972 7284 6978 7296
rect 7650 7284 7656 7296
rect 7708 7324 7714 7336
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 7708 7296 7757 7324
rect 7708 7284 7714 7296
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 9677 7327 9735 7333
rect 9677 7293 9689 7327
rect 9723 7324 9735 7327
rect 9723 7296 9996 7324
rect 9723 7293 9735 7296
rect 9677 7287 9735 7293
rect 9968 7200 9996 7296
rect 10042 7284 10048 7336
rect 10100 7324 10106 7336
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 10100 7296 10149 7324
rect 10100 7284 10106 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 10410 7284 10416 7336
rect 10468 7284 10474 7336
rect 10551 7327 10609 7333
rect 10551 7293 10563 7327
rect 10597 7324 10609 7327
rect 10870 7324 10876 7336
rect 10597 7296 10876 7324
rect 10597 7293 10609 7296
rect 10551 7287 10609 7293
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 11112 7296 11529 7324
rect 11112 7284 11118 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 13262 7284 13268 7336
rect 13320 7284 13326 7336
rect 2406 7148 2412 7200
rect 2464 7148 2470 7200
rect 9950 7148 9956 7200
rect 10008 7148 10014 7200
rect 10778 7148 10784 7200
rect 10836 7188 10842 7200
rect 11606 7188 11612 7200
rect 10836 7160 11612 7188
rect 10836 7148 10842 7160
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 1486 6944 1492 6996
rect 1544 6984 1550 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 1544 6956 2421 6984
rect 1544 6944 1550 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 3234 6944 3240 6996
rect 3292 6984 3298 6996
rect 8386 6984 8392 6996
rect 3292 6956 8392 6984
rect 3292 6944 3298 6956
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 10134 6944 10140 6996
rect 10192 6984 10198 6996
rect 11882 6984 11888 6996
rect 10192 6956 11888 6984
rect 10192 6944 10198 6956
rect 11882 6944 11888 6956
rect 11940 6984 11946 6996
rect 11940 6956 12296 6984
rect 11940 6944 11946 6956
rect 9398 6808 9404 6860
rect 9456 6808 9462 6860
rect 9858 6808 9864 6860
rect 9916 6808 9922 6860
rect 10134 6808 10140 6860
rect 10192 6808 10198 6860
rect 10318 6857 10324 6860
rect 10275 6851 10324 6857
rect 10275 6817 10287 6851
rect 10321 6817 10324 6851
rect 10275 6811 10324 6817
rect 10318 6808 10324 6811
rect 10376 6808 10382 6860
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 10594 6848 10600 6860
rect 10459 6820 10600 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 11701 6851 11759 6857
rect 11701 6817 11713 6851
rect 11747 6848 11759 6851
rect 12066 6848 12072 6860
rect 11747 6820 12072 6848
rect 11747 6817 11759 6820
rect 11701 6811 11759 6817
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 2314 6740 2320 6792
rect 2372 6740 2378 6792
rect 2406 6740 2412 6792
rect 2464 6780 2470 6792
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 2464 6752 2605 6780
rect 2464 6740 2470 6752
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 2593 6743 2651 6749
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 12268 6780 12296 6956
rect 13817 6919 13875 6925
rect 13817 6885 13829 6919
rect 13863 6885 13875 6919
rect 13817 6879 13875 6885
rect 13544 6860 13596 6866
rect 13832 6848 13860 6879
rect 15194 6848 15200 6860
rect 13832 6820 15200 6848
rect 15194 6808 15200 6820
rect 15252 6808 15258 6860
rect 13544 6802 13596 6808
rect 12805 6783 12863 6789
rect 12805 6780 12817 6783
rect 12268 6752 12817 6780
rect 11425 6743 11483 6749
rect 12805 6749 12817 6752
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 12943 6752 13492 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 1489 6715 1547 6721
rect 1489 6681 1501 6715
rect 1535 6712 1547 6715
rect 1535 6684 2176 6712
rect 1535 6681 1547 6684
rect 1489 6675 1547 6681
rect 842 6604 848 6656
rect 900 6644 906 6656
rect 2148 6653 2176 6684
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 900 6616 1593 6644
rect 900 6604 906 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6613 2191 6647
rect 9232 6644 9260 6740
rect 11440 6712 11468 6743
rect 12710 6712 12716 6724
rect 10888 6684 11284 6712
rect 11440 6684 12716 6712
rect 10888 6644 10916 6684
rect 9232 6616 10916 6644
rect 11057 6647 11115 6653
rect 2133 6607 2191 6613
rect 11057 6613 11069 6647
rect 11103 6644 11115 6647
rect 11146 6644 11152 6656
rect 11103 6616 11152 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 11256 6644 11284 6684
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 13265 6715 13323 6721
rect 13265 6681 13277 6715
rect 13311 6712 13323 6715
rect 13354 6712 13360 6724
rect 13311 6684 13360 6712
rect 13311 6681 13323 6684
rect 13265 6675 13323 6681
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 12526 6644 12532 6656
rect 11256 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 13464 6644 13492 6752
rect 13630 6672 13636 6724
rect 13688 6712 13694 6724
rect 14277 6715 14335 6721
rect 13688 6684 13952 6712
rect 13688 6672 13694 6684
rect 13814 6644 13820 6656
rect 13464 6616 13820 6644
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 13924 6644 13952 6684
rect 14277 6681 14289 6715
rect 14323 6712 14335 6715
rect 15102 6712 15108 6724
rect 14323 6684 15108 6712
rect 14323 6681 14335 6684
rect 14277 6675 14335 6681
rect 15102 6672 15108 6684
rect 15160 6672 15166 6724
rect 14369 6647 14427 6653
rect 14369 6644 14381 6647
rect 13924 6616 14381 6644
rect 14369 6613 14381 6616
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 2409 6443 2467 6449
rect 2409 6440 2421 6443
rect 2372 6412 2421 6440
rect 2372 6400 2378 6412
rect 2409 6409 2421 6412
rect 2455 6409 2467 6443
rect 2409 6403 2467 6409
rect 9125 6443 9183 6449
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 10042 6440 10048 6452
rect 9171 6412 10048 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11146 6400 11152 6452
rect 11204 6400 11210 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 14182 6440 14188 6452
rect 12768 6412 14188 6440
rect 12768 6400 12774 6412
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 11164 6372 11192 6400
rect 11164 6344 11560 6372
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 1578 6304 1584 6316
rect 1443 6276 1584 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 1671 6307 1729 6313
rect 1671 6273 1683 6307
rect 1717 6304 1729 6307
rect 5810 6304 5816 6316
rect 1717 6276 5816 6304
rect 1717 6273 1729 6276
rect 1671 6267 1729 6273
rect 5810 6264 5816 6276
rect 5868 6304 5874 6316
rect 8355 6307 8413 6313
rect 8355 6304 8367 6307
rect 5868 6276 8367 6304
rect 5868 6264 5874 6276
rect 8355 6273 8367 6276
rect 8401 6273 8413 6307
rect 8355 6267 8413 6273
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9088 6276 9505 6304
rect 9088 6264 9094 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 10686 6264 10692 6316
rect 10744 6264 10750 6316
rect 11532 6313 11560 6344
rect 13354 6332 13360 6384
rect 13412 6372 13418 6384
rect 14366 6372 14372 6384
rect 13412 6344 14372 6372
rect 13412 6332 13418 6344
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 12434 6264 12440 6316
rect 12492 6264 12498 6316
rect 12526 6264 12532 6316
rect 12584 6313 12590 6316
rect 12584 6307 12612 6313
rect 12600 6273 12612 6307
rect 12584 6267 12612 6273
rect 12584 6264 12590 6267
rect 12710 6264 12716 6316
rect 12768 6264 12774 6316
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7708 6208 8125 6236
rect 7708 6196 7714 6208
rect 8113 6205 8125 6208
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 9674 6196 9680 6248
rect 9732 6196 9738 6248
rect 9858 6196 9864 6248
rect 9916 6236 9922 6248
rect 10137 6239 10195 6245
rect 10137 6236 10149 6239
rect 9916 6208 10149 6236
rect 9916 6196 9922 6208
rect 10137 6205 10149 6208
rect 10183 6205 10195 6239
rect 10410 6236 10416 6248
rect 10137 6199 10195 6205
rect 10244 6208 10416 6236
rect 9692 6168 9720 6196
rect 9950 6168 9956 6180
rect 9692 6140 9956 6168
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 10244 6100 10272 6208
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10551 6239 10609 6245
rect 10551 6205 10563 6239
rect 10597 6236 10609 6239
rect 10870 6236 10876 6248
rect 10597 6208 10876 6236
rect 10597 6205 10609 6208
rect 10551 6199 10609 6205
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6236 11391 6239
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11379 6208 11713 6236
rect 11379 6205 11391 6208
rect 11333 6199 11391 6205
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 12158 6128 12164 6180
rect 12216 6128 12222 6180
rect 13372 6168 13400 6332
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6304 13691 6307
rect 14734 6304 14740 6316
rect 13679 6276 14740 6304
rect 13679 6273 13691 6276
rect 13633 6267 13691 6273
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 13906 6196 13912 6248
rect 13964 6196 13970 6248
rect 13096 6140 13400 6168
rect 13096 6100 13124 6140
rect 10244 6072 13124 6100
rect 13354 6060 13360 6112
rect 13412 6060 13418 6112
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 842 5856 848 5908
rect 900 5896 906 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 900 5868 1593 5896
rect 900 5856 906 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 8478 5856 8484 5908
rect 8536 5856 8542 5908
rect 9306 5856 9312 5908
rect 9364 5856 9370 5908
rect 11885 5899 11943 5905
rect 11885 5865 11897 5899
rect 11931 5896 11943 5899
rect 12710 5896 12716 5908
rect 11931 5868 12716 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 13262 5856 13268 5908
rect 13320 5856 13326 5908
rect 9324 5828 9352 5856
rect 8128 5800 9352 5828
rect 13909 5831 13967 5837
rect 4246 5760 4252 5772
rect 2056 5732 4252 5760
rect 2056 5701 2084 5732
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5692 2559 5695
rect 7469 5695 7527 5701
rect 2547 5664 2774 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5624 1547 5627
rect 2746 5624 2774 5664
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 7650 5692 7656 5704
rect 7515 5664 7656 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 7743 5695 7801 5701
rect 7743 5661 7755 5695
rect 7789 5692 7801 5695
rect 8128 5692 8156 5800
rect 13909 5797 13921 5831
rect 13955 5828 13967 5831
rect 14182 5828 14188 5840
rect 13955 5800 14188 5828
rect 13955 5797 13967 5800
rect 13909 5791 13967 5797
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 8202 5720 8208 5772
rect 8260 5760 8266 5772
rect 8260 5732 8432 5760
rect 8260 5720 8266 5732
rect 7789 5664 8156 5692
rect 7789 5661 7801 5664
rect 7743 5655 7801 5661
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8404 5692 8432 5732
rect 9766 5720 9772 5772
rect 9824 5760 9830 5772
rect 10778 5760 10784 5772
rect 9824 5732 10784 5760
rect 9824 5720 9830 5732
rect 10778 5720 10784 5732
rect 10836 5760 10842 5772
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 10836 5732 10885 5760
rect 10836 5720 10842 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 10873 5723 10931 5729
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12253 5763 12311 5769
rect 12253 5760 12265 5763
rect 12032 5732 12265 5760
rect 12032 5720 12038 5732
rect 12253 5729 12265 5732
rect 12299 5729 12311 5763
rect 12253 5723 12311 5729
rect 11115 5695 11173 5701
rect 11115 5692 11127 5695
rect 8404 5664 11127 5692
rect 11115 5661 11127 5664
rect 11161 5661 11173 5695
rect 11115 5655 11173 5661
rect 12495 5695 12553 5701
rect 12495 5661 12507 5695
rect 12541 5692 12553 5695
rect 12618 5692 12624 5704
rect 12541 5664 12624 5692
rect 12541 5661 12553 5664
rect 12495 5655 12553 5661
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 13354 5692 13360 5704
rect 13188 5664 13360 5692
rect 8312 5624 8340 5652
rect 1535 5596 2360 5624
rect 2746 5596 8340 5624
rect 1535 5593 1547 5596
rect 1489 5587 1547 5593
rect 2130 5516 2136 5568
rect 2188 5516 2194 5568
rect 2332 5565 2360 5596
rect 9306 5584 9312 5636
rect 9364 5624 9370 5636
rect 9364 5596 10088 5624
rect 9364 5584 9370 5596
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5525 2375 5559
rect 2317 5519 2375 5525
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 9950 5556 9956 5568
rect 4764 5528 9956 5556
rect 4764 5516 4770 5528
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10060 5556 10088 5596
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 13188 5624 13216 5664
rect 13354 5652 13360 5664
rect 13412 5692 13418 5704
rect 13998 5692 14004 5704
rect 13412 5664 14004 5692
rect 13412 5652 13418 5664
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 10928 5596 13216 5624
rect 10928 5584 10934 5596
rect 13722 5584 13728 5636
rect 13780 5584 13786 5636
rect 14277 5627 14335 5633
rect 14277 5593 14289 5627
rect 14323 5624 14335 5627
rect 15102 5624 15108 5636
rect 14323 5596 15108 5624
rect 14323 5593 14335 5596
rect 14277 5587 14335 5593
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 12802 5556 12808 5568
rect 10060 5528 12808 5556
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 14369 5559 14427 5565
rect 14369 5556 14381 5559
rect 13964 5528 14381 5556
rect 13964 5516 13970 5528
rect 14369 5525 14381 5528
rect 14415 5525 14427 5559
rect 14369 5519 14427 5525
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 9125 5355 9183 5361
rect 9125 5321 9137 5355
rect 9171 5352 9183 5355
rect 9858 5352 9864 5364
rect 9171 5324 9864 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 10505 5355 10563 5361
rect 10505 5321 10517 5355
rect 10551 5352 10563 5355
rect 10594 5352 10600 5364
rect 10551 5324 10600 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 13357 5355 13415 5361
rect 13357 5321 13369 5355
rect 13403 5352 13415 5355
rect 13538 5352 13544 5364
rect 13403 5324 13544 5352
rect 13403 5321 13415 5324
rect 13357 5315 13415 5321
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 1489 5287 1547 5293
rect 1489 5253 1501 5287
rect 1535 5284 1547 5287
rect 2130 5284 2136 5296
rect 1535 5256 2136 5284
rect 1535 5253 1547 5256
rect 1489 5247 1547 5253
rect 2130 5244 2136 5256
rect 2188 5244 2194 5296
rect 3602 5244 3608 5296
rect 3660 5284 3666 5296
rect 3660 5256 9720 5284
rect 3660 5244 3666 5256
rect 9692 5246 9720 5256
rect 7374 5176 7380 5228
rect 7432 5216 7438 5228
rect 7650 5216 7656 5228
rect 7432 5188 7656 5216
rect 7432 5176 7438 5188
rect 7650 5176 7656 5188
rect 7708 5216 7714 5228
rect 8113 5219 8171 5225
rect 8113 5216 8125 5219
rect 7708 5188 8125 5216
rect 7708 5176 7714 5188
rect 8113 5185 8125 5188
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 842 4972 848 5024
rect 900 5012 906 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 900 4984 1593 5012
rect 900 4972 906 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 8128 5012 8156 5179
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 9398 5216 9404 5228
rect 8444 5188 9404 5216
rect 8444 5176 8450 5188
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 9692 5225 9810 5246
rect 12619 5229 12677 5235
rect 9692 5219 9825 5225
rect 9692 5218 9779 5219
rect 9767 5185 9779 5218
rect 9813 5185 9825 5219
rect 9767 5179 9825 5185
rect 11974 5176 11980 5228
rect 12032 5216 12038 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 12032 5188 12357 5216
rect 12032 5176 12038 5188
rect 12345 5185 12357 5188
rect 12391 5216 12403 5219
rect 12526 5216 12532 5228
rect 12391 5188 12532 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 12619 5195 12631 5229
rect 12665 5216 12677 5229
rect 12710 5216 12716 5228
rect 12665 5195 12716 5216
rect 12619 5189 12716 5195
rect 12634 5188 12716 5189
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5117 9551 5151
rect 9493 5111 9551 5117
rect 9508 5012 9536 5111
rect 9766 5012 9772 5024
rect 8128 4984 9772 5012
rect 1581 4975 1639 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 3878 4808 3884 4820
rect 1627 4780 3884 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 11609 4811 11667 4817
rect 9456 4780 11284 4808
rect 9456 4768 9462 4780
rect 11256 4740 11284 4780
rect 11609 4777 11621 4811
rect 11655 4808 11667 4811
rect 12158 4808 12164 4820
rect 11655 4780 12164 4808
rect 11655 4777 11667 4780
rect 11609 4771 11667 4777
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 13446 4768 13452 4820
rect 13504 4808 13510 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13504 4780 13645 4808
rect 13504 4768 13510 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 11790 4740 11796 4752
rect 11256 4712 11796 4740
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 9916 4644 10609 4672
rect 9916 4632 9922 4644
rect 10597 4641 10609 4644
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 750 4564 756 4616
rect 808 4604 814 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 808 4576 1409 4604
rect 808 4564 814 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 10839 4607 10897 4613
rect 10839 4604 10851 4607
rect 1397 4567 1455 4573
rect 10704 4576 10851 4604
rect 8662 4496 8668 4548
rect 8720 4536 8726 4548
rect 10704 4536 10732 4576
rect 10839 4573 10851 4576
rect 10885 4573 10897 4607
rect 10839 4567 10897 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 12894 4613 12900 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 12584 4576 12633 4604
rect 12584 4564 12590 4576
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 12863 4607 12900 4613
rect 12863 4573 12875 4607
rect 12863 4567 12900 4573
rect 12894 4564 12900 4567
rect 12952 4564 12958 4616
rect 8720 4508 10732 4536
rect 8720 4496 8726 4508
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 13139 4131 13197 4137
rect 13139 4128 13151 4131
rect 11848 4100 13151 4128
rect 11848 4088 11854 4100
rect 13139 4097 13151 4100
rect 13185 4097 13197 4131
rect 13139 4091 13197 4097
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12584 4032 12909 4060
rect 12584 4020 12590 4032
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 13909 3927 13967 3933
rect 13909 3924 13921 3927
rect 13872 3896 13921 3924
rect 13872 3884 13878 3896
rect 13909 3893 13921 3896
rect 13955 3893 13967 3927
rect 13909 3887 13967 3893
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 9272 3692 14289 3720
rect 9272 3680 9278 3692
rect 14277 3689 14289 3692
rect 14323 3689 14335 3723
rect 14277 3683 14335 3689
rect 13354 3612 13360 3664
rect 13412 3612 13418 3664
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 12400 3556 13093 3584
rect 12400 3544 12406 3556
rect 13081 3553 13093 3556
rect 13127 3553 13139 3587
rect 13081 3547 13139 3553
rect 13372 3525 13400 3612
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3485 13415 3519
rect 13357 3479 13415 3485
rect 14182 3476 14188 3528
rect 14240 3476 14246 3528
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 13630 3000 13636 3052
rect 13688 3000 13694 3052
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3040 13967 3043
rect 14366 3040 14372 3052
rect 13955 3012 14372 3040
rect 13955 3009 13967 3012
rect 13909 3003 13967 3009
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
rect 5810 2048 5816 2100
rect 5868 2048 5874 2100
rect 6546 2048 6552 2100
rect 6604 2048 6610 2100
rect 7285 2091 7343 2097
rect 7285 2088 7297 2091
rect 6886 2060 7297 2088
rect 4062 1980 4068 2032
rect 4120 2020 4126 2032
rect 6886 2020 6914 2060
rect 7285 2057 7297 2060
rect 7331 2057 7343 2091
rect 7285 2051 7343 2057
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 8021 2091 8079 2097
rect 8021 2088 8033 2091
rect 7708 2060 8033 2088
rect 7708 2048 7714 2060
rect 8021 2057 8033 2060
rect 8067 2057 8079 2091
rect 8021 2051 8079 2057
rect 8846 2048 8852 2100
rect 8904 2088 8910 2100
rect 9401 2091 9459 2097
rect 9401 2088 9413 2091
rect 8904 2060 9413 2088
rect 8904 2048 8910 2060
rect 9401 2057 9413 2060
rect 9447 2057 9459 2091
rect 9401 2051 9459 2057
rect 9950 2048 9956 2100
rect 10008 2088 10014 2100
rect 10229 2091 10287 2097
rect 10229 2088 10241 2091
rect 10008 2060 10241 2088
rect 10008 2048 10014 2060
rect 10229 2057 10241 2060
rect 10275 2057 10287 2091
rect 10229 2051 10287 2057
rect 11701 2091 11759 2097
rect 11701 2057 11713 2091
rect 11747 2088 11759 2091
rect 11790 2088 11796 2100
rect 11747 2060 11796 2088
rect 11747 2057 11759 2060
rect 11701 2051 11759 2057
rect 11790 2048 11796 2060
rect 11848 2048 11854 2100
rect 12434 2048 12440 2100
rect 12492 2048 12498 2100
rect 14182 2048 14188 2100
rect 14240 2048 14246 2100
rect 4120 1992 6914 2020
rect 8757 2023 8815 2029
rect 4120 1980 4126 1992
rect 8757 1989 8769 2023
rect 8803 2020 8815 2023
rect 8938 2020 8944 2032
rect 8803 1992 8944 2020
rect 8803 1989 8815 1992
rect 8757 1983 8815 1989
rect 8938 1980 8944 1992
rect 8996 1980 9002 2032
rect 11054 1980 11060 2032
rect 11112 1980 11118 2032
rect 13446 1980 13452 2032
rect 13504 2020 13510 2032
rect 14093 2023 14151 2029
rect 14093 2020 14105 2023
rect 13504 1992 14105 2020
rect 13504 1980 13510 1992
rect 14093 1989 14105 1992
rect 14139 1989 14151 2023
rect 14093 1983 14151 1989
rect 1302 1912 1308 1964
rect 1360 1952 1366 1964
rect 1397 1955 1455 1961
rect 1397 1952 1409 1955
rect 1360 1924 1409 1952
rect 1360 1912 1366 1924
rect 1397 1921 1409 1924
rect 1443 1921 1455 1955
rect 1397 1915 1455 1921
rect 3050 1912 3056 1964
rect 3108 1912 3114 1964
rect 5718 1912 5724 1964
rect 5776 1912 5782 1964
rect 6454 1912 6460 1964
rect 6512 1912 6518 1964
rect 7190 1912 7196 1964
rect 7248 1912 7254 1964
rect 7926 1912 7932 1964
rect 7984 1912 7990 1964
rect 8570 1912 8576 1964
rect 8628 1912 8634 1964
rect 9306 1912 9312 1964
rect 9364 1912 9370 1964
rect 10134 1912 10140 1964
rect 10192 1912 10198 1964
rect 10870 1912 10876 1964
rect 10928 1912 10934 1964
rect 11606 1912 11612 1964
rect 11664 1912 11670 1964
rect 12342 1912 12348 1964
rect 12400 1912 12406 1964
rect 12989 1955 13047 1961
rect 12989 1921 13001 1955
rect 13035 1952 13047 1955
rect 13262 1952 13268 1964
rect 13035 1924 13268 1952
rect 13035 1921 13047 1924
rect 12989 1915 13047 1921
rect 13262 1912 13268 1924
rect 13320 1912 13326 1964
rect 13722 1912 13728 1964
rect 13780 1912 13786 1964
rect 2225 1887 2283 1893
rect 2225 1853 2237 1887
rect 2271 1853 2283 1887
rect 2225 1847 2283 1853
rect 3697 1887 3755 1893
rect 3697 1853 3709 1887
rect 3743 1884 3755 1887
rect 11146 1884 11152 1896
rect 3743 1856 11152 1884
rect 3743 1853 3755 1856
rect 3697 1847 3755 1853
rect 2240 1816 2268 1847
rect 11146 1844 11152 1856
rect 11204 1844 11210 1896
rect 13909 1887 13967 1893
rect 13909 1853 13921 1887
rect 13955 1884 13967 1887
rect 15194 1884 15200 1896
rect 13955 1856 15200 1884
rect 13955 1853 13967 1856
rect 13909 1847 13967 1853
rect 15194 1844 15200 1856
rect 15252 1844 15258 1896
rect 15378 1844 15384 1896
rect 15436 1844 15442 1896
rect 7374 1816 7380 1828
rect 2240 1788 7380 1816
rect 7374 1776 7380 1788
rect 7432 1776 7438 1828
rect 13173 1819 13231 1825
rect 13173 1785 13185 1819
rect 13219 1816 13231 1819
rect 15396 1816 15424 1844
rect 13219 1788 15424 1816
rect 13219 1785 13231 1788
rect 13173 1779 13231 1785
rect 1104 1658 14812 1680
rect 1104 1606 2663 1658
rect 2715 1606 2727 1658
rect 2779 1606 2791 1658
rect 2843 1606 2855 1658
rect 2907 1606 2919 1658
rect 2971 1606 6090 1658
rect 6142 1606 6154 1658
rect 6206 1606 6218 1658
rect 6270 1606 6282 1658
rect 6334 1606 6346 1658
rect 6398 1606 9517 1658
rect 9569 1606 9581 1658
rect 9633 1606 9645 1658
rect 9697 1606 9709 1658
rect 9761 1606 9773 1658
rect 9825 1606 12944 1658
rect 12996 1606 13008 1658
rect 13060 1606 13072 1658
rect 13124 1606 13136 1658
rect 13188 1606 13200 1658
rect 13252 1606 14812 1658
rect 1104 1584 14812 1606
rect 5718 1504 5724 1556
rect 5776 1544 5782 1556
rect 5813 1547 5871 1553
rect 5813 1544 5825 1547
rect 5776 1516 5825 1544
rect 5776 1504 5782 1516
rect 5813 1513 5825 1516
rect 5859 1513 5871 1547
rect 5813 1507 5871 1513
rect 6454 1504 6460 1556
rect 6512 1544 6518 1556
rect 6549 1547 6607 1553
rect 6549 1544 6561 1547
rect 6512 1516 6561 1544
rect 6512 1504 6518 1516
rect 6549 1513 6561 1516
rect 6595 1513 6607 1547
rect 6549 1507 6607 1513
rect 7190 1504 7196 1556
rect 7248 1544 7254 1556
rect 7285 1547 7343 1553
rect 7285 1544 7297 1547
rect 7248 1516 7297 1544
rect 7248 1504 7254 1516
rect 7285 1513 7297 1516
rect 7331 1513 7343 1547
rect 7285 1507 7343 1513
rect 7926 1504 7932 1556
rect 7984 1544 7990 1556
rect 8021 1547 8079 1553
rect 8021 1544 8033 1547
rect 7984 1516 8033 1544
rect 7984 1504 7990 1516
rect 8021 1513 8033 1516
rect 8067 1513 8079 1547
rect 8021 1507 8079 1513
rect 8570 1504 8576 1556
rect 8628 1544 8634 1556
rect 8941 1547 8999 1553
rect 8941 1544 8953 1547
rect 8628 1516 8953 1544
rect 8628 1504 8634 1516
rect 8941 1513 8953 1516
rect 8987 1513 8999 1547
rect 8941 1507 8999 1513
rect 9306 1504 9312 1556
rect 9364 1544 9370 1556
rect 9493 1547 9551 1553
rect 9493 1544 9505 1547
rect 9364 1516 9505 1544
rect 9364 1504 9370 1516
rect 9493 1513 9505 1516
rect 9539 1513 9551 1547
rect 9493 1507 9551 1513
rect 10134 1504 10140 1556
rect 10192 1544 10198 1556
rect 10229 1547 10287 1553
rect 10229 1544 10241 1547
rect 10192 1516 10241 1544
rect 10192 1504 10198 1516
rect 10229 1513 10241 1516
rect 10275 1513 10287 1547
rect 10229 1507 10287 1513
rect 10870 1504 10876 1556
rect 10928 1544 10934 1556
rect 10965 1547 11023 1553
rect 10965 1544 10977 1547
rect 10928 1516 10977 1544
rect 10928 1504 10934 1516
rect 10965 1513 10977 1516
rect 11011 1513 11023 1547
rect 10965 1507 11023 1513
rect 11606 1504 11612 1556
rect 11664 1544 11670 1556
rect 11701 1547 11759 1553
rect 11701 1544 11713 1547
rect 11664 1516 11713 1544
rect 11664 1504 11670 1516
rect 11701 1513 11713 1516
rect 11747 1513 11759 1547
rect 11701 1507 11759 1513
rect 12342 1504 12348 1556
rect 12400 1544 12406 1556
rect 12437 1547 12495 1553
rect 12437 1544 12449 1547
rect 12400 1516 12449 1544
rect 12400 1504 12406 1516
rect 12437 1513 12449 1516
rect 12483 1513 12495 1547
rect 12437 1507 12495 1513
rect 13173 1547 13231 1553
rect 13173 1513 13185 1547
rect 13219 1544 13231 1547
rect 13262 1544 13268 1556
rect 13219 1516 13268 1544
rect 13219 1513 13231 1516
rect 13173 1507 13231 1513
rect 13262 1504 13268 1516
rect 13320 1504 13326 1556
rect 13446 1504 13452 1556
rect 13504 1504 13510 1556
rect 13722 1504 13728 1556
rect 13780 1504 13786 1556
rect 12897 1479 12955 1485
rect 12897 1445 12909 1479
rect 12943 1445 12955 1479
rect 12897 1439 12955 1445
rect 2961 1411 3019 1417
rect 2961 1377 2973 1411
rect 3007 1408 3019 1411
rect 12526 1408 12532 1420
rect 3007 1380 12532 1408
rect 3007 1377 3019 1380
rect 2961 1371 3019 1377
rect 12526 1368 12532 1380
rect 12584 1368 12590 1420
rect 12912 1408 12940 1439
rect 12912 1380 13216 1408
rect 2130 1300 2136 1352
rect 2188 1300 2194 1352
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 4614 1300 4620 1352
rect 4672 1300 4678 1352
rect 5350 1300 5356 1352
rect 5408 1300 5414 1352
rect 5718 1300 5724 1352
rect 5776 1340 5782 1352
rect 5997 1343 6055 1349
rect 5997 1340 6009 1343
rect 5776 1312 6009 1340
rect 5776 1300 5782 1312
rect 5997 1309 6009 1312
rect 6043 1309 6055 1343
rect 5997 1303 6055 1309
rect 6454 1300 6460 1352
rect 6512 1340 6518 1352
rect 6733 1343 6791 1349
rect 6733 1340 6745 1343
rect 6512 1312 6745 1340
rect 6512 1300 6518 1312
rect 6733 1309 6745 1312
rect 6779 1309 6791 1343
rect 6733 1303 6791 1309
rect 7190 1300 7196 1352
rect 7248 1340 7254 1352
rect 7469 1343 7527 1349
rect 7469 1340 7481 1343
rect 7248 1312 7481 1340
rect 7248 1300 7254 1312
rect 7469 1309 7481 1312
rect 7515 1309 7527 1343
rect 7469 1303 7527 1309
rect 8202 1300 8208 1352
rect 8260 1300 8266 1352
rect 8662 1300 8668 1352
rect 8720 1340 8726 1352
rect 9125 1343 9183 1349
rect 9125 1340 9137 1343
rect 8720 1312 9137 1340
rect 8720 1300 8726 1312
rect 9125 1309 9137 1312
rect 9171 1309 9183 1343
rect 9125 1303 9183 1309
rect 9674 1300 9680 1352
rect 9732 1300 9738 1352
rect 10134 1300 10140 1352
rect 10192 1340 10198 1352
rect 10413 1343 10471 1349
rect 10413 1340 10425 1343
rect 10192 1312 10425 1340
rect 10192 1300 10198 1312
rect 10413 1309 10425 1312
rect 10459 1309 10471 1343
rect 10413 1303 10471 1309
rect 10870 1300 10876 1352
rect 10928 1340 10934 1352
rect 11149 1343 11207 1349
rect 11149 1340 11161 1343
rect 10928 1312 11161 1340
rect 10928 1300 10934 1312
rect 11149 1309 11161 1312
rect 11195 1309 11207 1343
rect 11149 1303 11207 1309
rect 11606 1300 11612 1352
rect 11664 1340 11670 1352
rect 11885 1343 11943 1349
rect 11885 1340 11897 1343
rect 11664 1312 11897 1340
rect 11664 1300 11670 1312
rect 11885 1309 11897 1312
rect 11931 1309 11943 1343
rect 11885 1303 11943 1309
rect 12342 1300 12348 1352
rect 12400 1340 12406 1352
rect 12621 1343 12679 1349
rect 12621 1340 12633 1343
rect 12400 1312 12633 1340
rect 12400 1300 12406 1312
rect 12621 1309 12633 1312
rect 12667 1309 12679 1343
rect 12621 1303 12679 1309
rect 13081 1343 13139 1349
rect 13081 1309 13093 1343
rect 13127 1309 13139 1343
rect 13081 1303 13139 1309
rect 1578 1232 1584 1284
rect 1636 1272 1642 1284
rect 4065 1275 4123 1281
rect 4065 1272 4077 1275
rect 1636 1244 4077 1272
rect 1636 1232 1642 1244
rect 4065 1241 4077 1244
rect 4111 1241 4123 1275
rect 4065 1235 4123 1241
rect 4246 1232 4252 1284
rect 4304 1272 4310 1284
rect 4433 1275 4491 1281
rect 4433 1272 4445 1275
rect 4304 1244 4445 1272
rect 4304 1232 4310 1244
rect 4433 1241 4445 1244
rect 4479 1241 4491 1275
rect 4433 1235 4491 1241
rect 5166 1232 5172 1284
rect 5224 1232 5230 1284
rect 13096 1204 13124 1303
rect 13188 1272 13216 1380
rect 13832 1380 14044 1408
rect 13354 1300 13360 1352
rect 13412 1300 13418 1352
rect 13633 1343 13691 1349
rect 13633 1309 13645 1343
rect 13679 1340 13691 1343
rect 13832 1340 13860 1380
rect 13679 1312 13860 1340
rect 13679 1309 13691 1312
rect 13633 1303 13691 1309
rect 13906 1300 13912 1352
rect 13964 1300 13970 1352
rect 14016 1340 14044 1380
rect 14550 1340 14556 1352
rect 14016 1312 14556 1340
rect 14550 1300 14556 1312
rect 14608 1300 14614 1352
rect 15286 1300 15292 1352
rect 15344 1300 15350 1352
rect 14185 1275 14243 1281
rect 14185 1272 14197 1275
rect 13188 1244 14197 1272
rect 14185 1241 14197 1244
rect 14231 1241 14243 1275
rect 14185 1235 14243 1241
rect 14369 1275 14427 1281
rect 14369 1241 14381 1275
rect 14415 1272 14427 1275
rect 15304 1272 15332 1300
rect 14415 1244 15332 1272
rect 14415 1241 14427 1244
rect 14369 1235 14427 1241
rect 15286 1204 15292 1216
rect 13096 1176 15292 1204
rect 15286 1164 15292 1176
rect 15344 1164 15350 1216
rect 1104 1114 14971 1136
rect 1104 1062 4376 1114
rect 4428 1062 4440 1114
rect 4492 1062 4504 1114
rect 4556 1062 4568 1114
rect 4620 1062 4632 1114
rect 4684 1062 7803 1114
rect 7855 1062 7867 1114
rect 7919 1062 7931 1114
rect 7983 1062 7995 1114
rect 8047 1062 8059 1114
rect 8111 1062 11230 1114
rect 11282 1062 11294 1114
rect 11346 1062 11358 1114
rect 11410 1062 11422 1114
rect 11474 1062 11486 1114
rect 11538 1062 14657 1114
rect 14709 1062 14721 1114
rect 14773 1062 14785 1114
rect 14837 1062 14849 1114
rect 14901 1062 14913 1114
rect 14965 1062 14971 1114
rect 1104 1040 14971 1062
<< via1 >>
rect 4376 43494 4428 43546
rect 4440 43494 4492 43546
rect 4504 43494 4556 43546
rect 4568 43494 4620 43546
rect 4632 43494 4684 43546
rect 7803 43494 7855 43546
rect 7867 43494 7919 43546
rect 7931 43494 7983 43546
rect 7995 43494 8047 43546
rect 8059 43494 8111 43546
rect 11230 43494 11282 43546
rect 11294 43494 11346 43546
rect 11358 43494 11410 43546
rect 11422 43494 11474 43546
rect 11486 43494 11538 43546
rect 14657 43494 14709 43546
rect 14721 43494 14773 43546
rect 14785 43494 14837 43546
rect 14849 43494 14901 43546
rect 14913 43494 14965 43546
rect 1584 43435 1636 43444
rect 1584 43401 1593 43435
rect 1593 43401 1627 43435
rect 1627 43401 1636 43435
rect 1584 43392 1636 43401
rect 2320 43435 2372 43444
rect 2320 43401 2329 43435
rect 2329 43401 2363 43435
rect 2363 43401 2372 43435
rect 2320 43392 2372 43401
rect 2872 43435 2924 43444
rect 2872 43401 2881 43435
rect 2881 43401 2915 43435
rect 2915 43401 2924 43435
rect 2872 43392 2924 43401
rect 848 43324 900 43376
rect 3516 43392 3568 43444
rect 4252 43392 4304 43444
rect 5264 43435 5316 43444
rect 5264 43401 5273 43435
rect 5273 43401 5307 43435
rect 5307 43401 5316 43435
rect 5264 43392 5316 43401
rect 5908 43435 5960 43444
rect 5908 43401 5917 43435
rect 5917 43401 5951 43435
rect 5951 43401 5960 43435
rect 5908 43392 5960 43401
rect 6736 43435 6788 43444
rect 6736 43401 6745 43435
rect 6745 43401 6779 43435
rect 6779 43401 6788 43435
rect 6736 43392 6788 43401
rect 7472 43435 7524 43444
rect 7472 43401 7481 43435
rect 7481 43401 7515 43435
rect 7515 43401 7524 43435
rect 7472 43392 7524 43401
rect 8208 43435 8260 43444
rect 8208 43401 8217 43435
rect 8217 43401 8251 43435
rect 8251 43401 8260 43435
rect 8208 43392 8260 43401
rect 8668 43392 8720 43444
rect 9404 43392 9456 43444
rect 10416 43435 10468 43444
rect 10416 43401 10425 43435
rect 10425 43401 10459 43435
rect 10459 43401 10468 43435
rect 10416 43392 10468 43401
rect 10876 43392 10928 43444
rect 11888 43392 11940 43444
rect 12348 43392 12400 43444
rect 13084 43392 13136 43444
rect 15292 43392 15344 43444
rect 1768 43256 1820 43308
rect 2136 43299 2188 43308
rect 2136 43265 2145 43299
rect 2145 43265 2179 43299
rect 2179 43265 2188 43299
rect 2136 43256 2188 43265
rect 3056 43256 3108 43308
rect 3240 43299 3292 43308
rect 3240 43265 3249 43299
rect 3249 43265 3283 43299
rect 3283 43265 3292 43299
rect 3240 43256 3292 43265
rect 3792 43299 3844 43308
rect 3792 43265 3801 43299
rect 3801 43265 3835 43299
rect 3835 43265 3844 43299
rect 3792 43256 3844 43265
rect 4436 43299 4488 43308
rect 4436 43265 4445 43299
rect 4445 43265 4479 43299
rect 4479 43265 4488 43299
rect 4436 43256 4488 43265
rect 5080 43299 5132 43308
rect 5080 43265 5089 43299
rect 5089 43265 5123 43299
rect 5123 43265 5132 43299
rect 5080 43256 5132 43265
rect 5816 43299 5868 43308
rect 5816 43265 5825 43299
rect 5825 43265 5859 43299
rect 5859 43265 5868 43299
rect 5816 43256 5868 43265
rect 6644 43299 6696 43308
rect 6644 43265 6653 43299
rect 6653 43265 6687 43299
rect 6687 43265 6696 43299
rect 6644 43256 6696 43265
rect 7288 43299 7340 43308
rect 7288 43265 7297 43299
rect 7297 43265 7331 43299
rect 7331 43265 7340 43299
rect 7288 43256 7340 43265
rect 8116 43299 8168 43308
rect 8116 43265 8125 43299
rect 8125 43265 8159 43299
rect 8159 43265 8168 43299
rect 8116 43256 8168 43265
rect 8944 43299 8996 43308
rect 8944 43265 8953 43299
rect 8953 43265 8987 43299
rect 8987 43265 8996 43299
rect 8944 43256 8996 43265
rect 9220 43256 9272 43308
rect 10232 43299 10284 43308
rect 10232 43265 10241 43299
rect 10241 43265 10275 43299
rect 10275 43265 10284 43299
rect 10232 43256 10284 43265
rect 11612 43299 11664 43308
rect 11612 43265 11621 43299
rect 11621 43265 11655 43299
rect 11655 43265 11664 43299
rect 11612 43256 11664 43265
rect 12072 43299 12124 43308
rect 12072 43265 12081 43299
rect 12081 43265 12115 43299
rect 12115 43265 12124 43299
rect 12072 43256 12124 43265
rect 12532 43299 12584 43308
rect 12532 43265 12541 43299
rect 12541 43265 12575 43299
rect 12575 43265 12584 43299
rect 12532 43256 12584 43265
rect 12808 43256 12860 43308
rect 13728 43256 13780 43308
rect 15016 43256 15068 43308
rect 14096 43095 14148 43104
rect 14096 43061 14105 43095
rect 14105 43061 14139 43095
rect 14139 43061 14148 43095
rect 14096 43052 14148 43061
rect 2663 42950 2715 43002
rect 2727 42950 2779 43002
rect 2791 42950 2843 43002
rect 2855 42950 2907 43002
rect 2919 42950 2971 43002
rect 6090 42950 6142 43002
rect 6154 42950 6206 43002
rect 6218 42950 6270 43002
rect 6282 42950 6334 43002
rect 6346 42950 6398 43002
rect 9517 42950 9569 43002
rect 9581 42950 9633 43002
rect 9645 42950 9697 43002
rect 9709 42950 9761 43002
rect 9773 42950 9825 43002
rect 12944 42950 12996 43002
rect 13008 42950 13060 43002
rect 13072 42950 13124 43002
rect 13136 42950 13188 43002
rect 13200 42950 13252 43002
rect 3240 42848 3292 42900
rect 3792 42848 3844 42900
rect 4436 42848 4488 42900
rect 5080 42848 5132 42900
rect 5816 42848 5868 42900
rect 6644 42848 6696 42900
rect 7288 42848 7340 42900
rect 8116 42848 8168 42900
rect 8944 42848 8996 42900
rect 9220 42891 9272 42900
rect 9220 42857 9229 42891
rect 9229 42857 9263 42891
rect 9263 42857 9272 42891
rect 9220 42848 9272 42857
rect 10232 42891 10284 42900
rect 10232 42857 10241 42891
rect 10241 42857 10275 42891
rect 10275 42857 10284 42891
rect 10232 42848 10284 42857
rect 11612 42848 11664 42900
rect 12072 42848 12124 42900
rect 12532 42848 12584 42900
rect 12808 42848 12860 42900
rect 3792 42712 3844 42764
rect 3516 42687 3568 42696
rect 3516 42653 3525 42687
rect 3525 42653 3559 42687
rect 3559 42653 3568 42687
rect 3516 42644 3568 42653
rect 4068 42644 4120 42696
rect 5080 42687 5132 42696
rect 5080 42653 5089 42687
rect 5089 42653 5123 42687
rect 5123 42653 5132 42687
rect 5080 42644 5132 42653
rect 14556 42712 14608 42764
rect 4804 42576 4856 42628
rect 3976 42508 4028 42560
rect 7288 42687 7340 42696
rect 7288 42653 7297 42687
rect 7297 42653 7331 42687
rect 7331 42653 7340 42687
rect 7288 42644 7340 42653
rect 7472 42644 7524 42696
rect 7196 42576 7248 42628
rect 9404 42687 9456 42696
rect 9404 42653 9413 42687
rect 9413 42653 9447 42687
rect 9447 42653 9456 42687
rect 9404 42644 9456 42653
rect 8852 42508 8904 42560
rect 10968 42687 11020 42696
rect 10968 42653 10977 42687
rect 10977 42653 11011 42687
rect 11011 42653 11020 42687
rect 10968 42644 11020 42653
rect 11704 42687 11756 42696
rect 11704 42653 11713 42687
rect 11713 42653 11747 42687
rect 11747 42653 11756 42687
rect 11704 42644 11756 42653
rect 12440 42687 12492 42696
rect 12440 42653 12449 42687
rect 12449 42653 12483 42687
rect 12483 42653 12492 42687
rect 12440 42644 12492 42653
rect 13544 42619 13596 42628
rect 13544 42585 13553 42619
rect 13553 42585 13587 42619
rect 13587 42585 13596 42619
rect 13544 42576 13596 42585
rect 15292 42644 15344 42696
rect 15200 42576 15252 42628
rect 13728 42508 13780 42560
rect 4376 42406 4428 42458
rect 4440 42406 4492 42458
rect 4504 42406 4556 42458
rect 4568 42406 4620 42458
rect 4632 42406 4684 42458
rect 7803 42406 7855 42458
rect 7867 42406 7919 42458
rect 7931 42406 7983 42458
rect 7995 42406 8047 42458
rect 8059 42406 8111 42458
rect 11230 42406 11282 42458
rect 11294 42406 11346 42458
rect 11358 42406 11410 42458
rect 11422 42406 11474 42458
rect 11486 42406 11538 42458
rect 14657 42406 14709 42458
rect 14721 42406 14773 42458
rect 14785 42406 14837 42458
rect 14849 42406 14901 42458
rect 14913 42406 14965 42458
rect 2136 42304 2188 42356
rect 4068 42347 4120 42356
rect 4068 42313 4077 42347
rect 4077 42313 4111 42347
rect 4111 42313 4120 42347
rect 4068 42304 4120 42313
rect 5080 42304 5132 42356
rect 3884 42236 3936 42288
rect 7196 42304 7248 42356
rect 7288 42304 7340 42356
rect 7472 42304 7524 42356
rect 13544 42304 13596 42356
rect 13820 42304 13872 42356
rect 2228 42211 2280 42220
rect 2228 42177 2237 42211
rect 2237 42177 2271 42211
rect 2271 42177 2280 42211
rect 2228 42168 2280 42177
rect 4252 42211 4304 42220
rect 4252 42177 4261 42211
rect 4261 42177 4295 42211
rect 4295 42177 4304 42211
rect 4252 42168 4304 42177
rect 5080 42211 5132 42220
rect 5080 42177 5089 42211
rect 5089 42177 5123 42211
rect 5123 42177 5132 42211
rect 5080 42168 5132 42177
rect 4068 42100 4120 42152
rect 1032 42032 1084 42084
rect 14096 42279 14148 42288
rect 14096 42245 14105 42279
rect 14105 42245 14139 42279
rect 14139 42245 14148 42279
rect 14096 42236 14148 42245
rect 13912 42211 13964 42220
rect 13912 42177 13921 42211
rect 13921 42177 13955 42211
rect 13955 42177 13964 42211
rect 13912 42168 13964 42177
rect 2663 41862 2715 41914
rect 2727 41862 2779 41914
rect 2791 41862 2843 41914
rect 2855 41862 2907 41914
rect 2919 41862 2971 41914
rect 6090 41862 6142 41914
rect 6154 41862 6206 41914
rect 6218 41862 6270 41914
rect 6282 41862 6334 41914
rect 6346 41862 6398 41914
rect 9517 41862 9569 41914
rect 9581 41862 9633 41914
rect 9645 41862 9697 41914
rect 9709 41862 9761 41914
rect 9773 41862 9825 41914
rect 12944 41862 12996 41914
rect 13008 41862 13060 41914
rect 13072 41862 13124 41914
rect 13136 41862 13188 41914
rect 13200 41862 13252 41914
rect 4160 41760 4212 41812
rect 8852 41760 8904 41812
rect 4376 41318 4428 41370
rect 4440 41318 4492 41370
rect 4504 41318 4556 41370
rect 4568 41318 4620 41370
rect 4632 41318 4684 41370
rect 7803 41318 7855 41370
rect 7867 41318 7919 41370
rect 7931 41318 7983 41370
rect 7995 41318 8047 41370
rect 8059 41318 8111 41370
rect 11230 41318 11282 41370
rect 11294 41318 11346 41370
rect 11358 41318 11410 41370
rect 11422 41318 11474 41370
rect 11486 41318 11538 41370
rect 14657 41318 14709 41370
rect 14721 41318 14773 41370
rect 14785 41318 14837 41370
rect 14849 41318 14901 41370
rect 14913 41318 14965 41370
rect 756 41080 808 41132
rect 9312 40876 9364 40928
rect 2663 40774 2715 40826
rect 2727 40774 2779 40826
rect 2791 40774 2843 40826
rect 2855 40774 2907 40826
rect 2919 40774 2971 40826
rect 6090 40774 6142 40826
rect 6154 40774 6206 40826
rect 6218 40774 6270 40826
rect 6282 40774 6334 40826
rect 6346 40774 6398 40826
rect 9517 40774 9569 40826
rect 9581 40774 9633 40826
rect 9645 40774 9697 40826
rect 9709 40774 9761 40826
rect 9773 40774 9825 40826
rect 12944 40774 12996 40826
rect 13008 40774 13060 40826
rect 13072 40774 13124 40826
rect 13136 40774 13188 40826
rect 13200 40774 13252 40826
rect 756 40468 808 40520
rect 13544 40443 13596 40452
rect 13544 40409 13553 40443
rect 13553 40409 13587 40443
rect 13587 40409 13596 40443
rect 13544 40400 13596 40409
rect 5172 40332 5224 40384
rect 13728 40332 13780 40384
rect 4376 40230 4428 40282
rect 4440 40230 4492 40282
rect 4504 40230 4556 40282
rect 4568 40230 4620 40282
rect 4632 40230 4684 40282
rect 7803 40230 7855 40282
rect 7867 40230 7919 40282
rect 7931 40230 7983 40282
rect 7995 40230 8047 40282
rect 8059 40230 8111 40282
rect 11230 40230 11282 40282
rect 11294 40230 11346 40282
rect 11358 40230 11410 40282
rect 11422 40230 11474 40282
rect 11486 40230 11538 40282
rect 14657 40230 14709 40282
rect 14721 40230 14773 40282
rect 14785 40230 14837 40282
rect 14849 40230 14901 40282
rect 14913 40230 14965 40282
rect 13544 40128 13596 40180
rect 9312 39992 9364 40044
rect 13360 40035 13412 40044
rect 13360 40001 13369 40035
rect 13369 40001 13403 40035
rect 13403 40001 13412 40035
rect 13360 39992 13412 40001
rect 13912 40035 13964 40044
rect 13912 40001 13921 40035
rect 13921 40001 13955 40035
rect 13955 40001 13964 40035
rect 13912 39992 13964 40001
rect 14004 39788 14056 39840
rect 14188 39831 14240 39840
rect 14188 39797 14197 39831
rect 14197 39797 14231 39831
rect 14231 39797 14240 39831
rect 14188 39788 14240 39797
rect 2663 39686 2715 39738
rect 2727 39686 2779 39738
rect 2791 39686 2843 39738
rect 2855 39686 2907 39738
rect 2919 39686 2971 39738
rect 6090 39686 6142 39738
rect 6154 39686 6206 39738
rect 6218 39686 6270 39738
rect 6282 39686 6334 39738
rect 6346 39686 6398 39738
rect 9517 39686 9569 39738
rect 9581 39686 9633 39738
rect 9645 39686 9697 39738
rect 9709 39686 9761 39738
rect 9773 39686 9825 39738
rect 12944 39686 12996 39738
rect 13008 39686 13060 39738
rect 13072 39686 13124 39738
rect 13136 39686 13188 39738
rect 13200 39686 13252 39738
rect 13360 39584 13412 39636
rect 13912 39516 13964 39568
rect 756 39380 808 39432
rect 5172 39380 5224 39432
rect 12808 39380 12860 39432
rect 13268 39380 13320 39432
rect 1584 39287 1636 39296
rect 1584 39253 1593 39287
rect 1593 39253 1627 39287
rect 1627 39253 1636 39287
rect 1584 39244 1636 39253
rect 13544 39355 13596 39364
rect 13544 39321 13553 39355
rect 13553 39321 13587 39355
rect 13587 39321 13596 39355
rect 13544 39312 13596 39321
rect 13912 39355 13964 39364
rect 13912 39321 13921 39355
rect 13921 39321 13955 39355
rect 13955 39321 13964 39355
rect 13912 39312 13964 39321
rect 14372 39287 14424 39296
rect 14372 39253 14381 39287
rect 14381 39253 14415 39287
rect 14415 39253 14424 39287
rect 14372 39244 14424 39253
rect 4376 39142 4428 39194
rect 4440 39142 4492 39194
rect 4504 39142 4556 39194
rect 4568 39142 4620 39194
rect 4632 39142 4684 39194
rect 7803 39142 7855 39194
rect 7867 39142 7919 39194
rect 7931 39142 7983 39194
rect 7995 39142 8047 39194
rect 8059 39142 8111 39194
rect 11230 39142 11282 39194
rect 11294 39142 11346 39194
rect 11358 39142 11410 39194
rect 11422 39142 11474 39194
rect 11486 39142 11538 39194
rect 14657 39142 14709 39194
rect 14721 39142 14773 39194
rect 14785 39142 14837 39194
rect 14849 39142 14901 39194
rect 14913 39142 14965 39194
rect 1584 39040 1636 39092
rect 13544 39040 13596 39092
rect 12808 38972 12860 39024
rect 1400 38947 1452 38956
rect 1400 38913 1409 38947
rect 1409 38913 1443 38947
rect 1443 38913 1452 38947
rect 1400 38904 1452 38913
rect 12716 38904 12768 38956
rect 12348 38836 12400 38888
rect 13360 38947 13412 38956
rect 13360 38913 13369 38947
rect 13369 38913 13403 38947
rect 13403 38913 13412 38947
rect 13360 38904 13412 38913
rect 14004 38904 14056 38956
rect 13544 38836 13596 38888
rect 13820 38768 13872 38820
rect 12808 38700 12860 38752
rect 13636 38743 13688 38752
rect 13636 38709 13645 38743
rect 13645 38709 13679 38743
rect 13679 38709 13688 38743
rect 13636 38700 13688 38709
rect 14188 38743 14240 38752
rect 14188 38709 14197 38743
rect 14197 38709 14231 38743
rect 14231 38709 14240 38743
rect 14188 38700 14240 38709
rect 2663 38598 2715 38650
rect 2727 38598 2779 38650
rect 2791 38598 2843 38650
rect 2855 38598 2907 38650
rect 2919 38598 2971 38650
rect 6090 38598 6142 38650
rect 6154 38598 6206 38650
rect 6218 38598 6270 38650
rect 6282 38598 6334 38650
rect 6346 38598 6398 38650
rect 9517 38598 9569 38650
rect 9581 38598 9633 38650
rect 9645 38598 9697 38650
rect 9709 38598 9761 38650
rect 9773 38598 9825 38650
rect 12944 38598 12996 38650
rect 13008 38598 13060 38650
rect 13072 38598 13124 38650
rect 13136 38598 13188 38650
rect 13200 38598 13252 38650
rect 12716 38539 12768 38548
rect 12716 38505 12725 38539
rect 12725 38505 12759 38539
rect 12759 38505 12768 38539
rect 12716 38496 12768 38505
rect 13268 38496 13320 38548
rect 12716 38360 12768 38412
rect 12624 38335 12676 38344
rect 12624 38301 12633 38335
rect 12633 38301 12667 38335
rect 12667 38301 12676 38335
rect 12624 38292 12676 38301
rect 13452 38335 13504 38344
rect 13452 38301 13461 38335
rect 13461 38301 13495 38335
rect 13495 38301 13504 38335
rect 13452 38292 13504 38301
rect 13820 38292 13872 38344
rect 12808 38156 12860 38208
rect 13268 38199 13320 38208
rect 13268 38165 13277 38199
rect 13277 38165 13311 38199
rect 13311 38165 13320 38199
rect 13268 38156 13320 38165
rect 13820 38199 13872 38208
rect 13820 38165 13829 38199
rect 13829 38165 13863 38199
rect 13863 38165 13872 38199
rect 13820 38156 13872 38165
rect 14372 38199 14424 38208
rect 14372 38165 14381 38199
rect 14381 38165 14415 38199
rect 14415 38165 14424 38199
rect 14372 38156 14424 38165
rect 4376 38054 4428 38106
rect 4440 38054 4492 38106
rect 4504 38054 4556 38106
rect 4568 38054 4620 38106
rect 4632 38054 4684 38106
rect 7803 38054 7855 38106
rect 7867 38054 7919 38106
rect 7931 38054 7983 38106
rect 7995 38054 8047 38106
rect 8059 38054 8111 38106
rect 11230 38054 11282 38106
rect 11294 38054 11346 38106
rect 11358 38054 11410 38106
rect 11422 38054 11474 38106
rect 11486 38054 11538 38106
rect 14657 38054 14709 38106
rect 14721 38054 14773 38106
rect 14785 38054 14837 38106
rect 14849 38054 14901 38106
rect 14913 38054 14965 38106
rect 12624 37952 12676 38004
rect 756 37816 808 37868
rect 10784 37816 10836 37868
rect 13268 37884 13320 37936
rect 14004 37884 14056 37936
rect 7656 37680 7708 37732
rect 12624 37748 12676 37800
rect 13544 37859 13596 37868
rect 13544 37825 13553 37859
rect 13553 37825 13587 37859
rect 13587 37825 13596 37859
rect 13544 37816 13596 37825
rect 14004 37748 14056 37800
rect 12256 37680 12308 37732
rect 13360 37612 13412 37664
rect 13728 37612 13780 37664
rect 15108 37612 15160 37664
rect 2663 37510 2715 37562
rect 2727 37510 2779 37562
rect 2791 37510 2843 37562
rect 2855 37510 2907 37562
rect 2919 37510 2971 37562
rect 6090 37510 6142 37562
rect 6154 37510 6206 37562
rect 6218 37510 6270 37562
rect 6282 37510 6334 37562
rect 6346 37510 6398 37562
rect 9517 37510 9569 37562
rect 9581 37510 9633 37562
rect 9645 37510 9697 37562
rect 9709 37510 9761 37562
rect 9773 37510 9825 37562
rect 12944 37510 12996 37562
rect 13008 37510 13060 37562
rect 13072 37510 13124 37562
rect 13136 37510 13188 37562
rect 13200 37510 13252 37562
rect 10784 37451 10836 37460
rect 10784 37417 10793 37451
rect 10793 37417 10827 37451
rect 10827 37417 10836 37451
rect 10784 37408 10836 37417
rect 12624 37451 12676 37460
rect 12624 37417 12633 37451
rect 12633 37417 12667 37451
rect 12667 37417 12676 37451
rect 12624 37408 12676 37417
rect 13544 37408 13596 37460
rect 10508 37272 10560 37324
rect 12532 37247 12584 37256
rect 12532 37213 12541 37247
rect 12541 37213 12575 37247
rect 12575 37213 12584 37247
rect 12532 37204 12584 37213
rect 15384 37272 15436 37324
rect 13084 37247 13136 37256
rect 13084 37213 13093 37247
rect 13093 37213 13127 37247
rect 13127 37213 13136 37247
rect 13084 37204 13136 37213
rect 13360 37247 13412 37256
rect 13360 37213 13369 37247
rect 13369 37213 13403 37247
rect 13403 37213 13412 37247
rect 13360 37204 13412 37213
rect 756 37136 808 37188
rect 9128 37136 9180 37188
rect 12348 37111 12400 37120
rect 12348 37077 12357 37111
rect 12357 37077 12391 37111
rect 12391 37077 12400 37111
rect 12348 37068 12400 37077
rect 13084 37068 13136 37120
rect 14372 37111 14424 37120
rect 14372 37077 14381 37111
rect 14381 37077 14415 37111
rect 14415 37077 14424 37111
rect 14372 37068 14424 37077
rect 4376 36966 4428 37018
rect 4440 36966 4492 37018
rect 4504 36966 4556 37018
rect 4568 36966 4620 37018
rect 4632 36966 4684 37018
rect 7803 36966 7855 37018
rect 7867 36966 7919 37018
rect 7931 36966 7983 37018
rect 7995 36966 8047 37018
rect 8059 36966 8111 37018
rect 11230 36966 11282 37018
rect 11294 36966 11346 37018
rect 11358 36966 11410 37018
rect 11422 36966 11474 37018
rect 11486 36966 11538 37018
rect 14657 36966 14709 37018
rect 14721 36966 14773 37018
rect 14785 36966 14837 37018
rect 14849 36966 14901 37018
rect 14913 36966 14965 37018
rect 12624 36864 12676 36916
rect 13084 36864 13136 36916
rect 11060 36728 11112 36780
rect 12164 36728 12216 36780
rect 10140 36660 10192 36712
rect 12716 36728 12768 36780
rect 13636 36796 13688 36848
rect 13820 36728 13872 36780
rect 14004 36728 14056 36780
rect 12256 36592 12308 36644
rect 12348 36592 12400 36644
rect 13268 36660 13320 36712
rect 12440 36567 12492 36576
rect 12440 36533 12449 36567
rect 12449 36533 12483 36567
rect 12483 36533 12492 36567
rect 12440 36524 12492 36533
rect 13728 36567 13780 36576
rect 13728 36533 13737 36567
rect 13737 36533 13771 36567
rect 13771 36533 13780 36567
rect 13728 36524 13780 36533
rect 2663 36422 2715 36474
rect 2727 36422 2779 36474
rect 2791 36422 2843 36474
rect 2855 36422 2907 36474
rect 2919 36422 2971 36474
rect 6090 36422 6142 36474
rect 6154 36422 6206 36474
rect 6218 36422 6270 36474
rect 6282 36422 6334 36474
rect 6346 36422 6398 36474
rect 9517 36422 9569 36474
rect 9581 36422 9633 36474
rect 9645 36422 9697 36474
rect 9709 36422 9761 36474
rect 9773 36422 9825 36474
rect 12944 36422 12996 36474
rect 13008 36422 13060 36474
rect 13072 36422 13124 36474
rect 13136 36422 13188 36474
rect 13200 36422 13252 36474
rect 9128 36363 9180 36372
rect 9128 36329 9137 36363
rect 9137 36329 9171 36363
rect 9171 36329 9180 36363
rect 9128 36320 9180 36329
rect 12164 36320 12216 36372
rect 12348 36363 12400 36372
rect 12348 36329 12357 36363
rect 12357 36329 12391 36363
rect 12391 36329 12400 36363
rect 12348 36320 12400 36329
rect 12716 36320 12768 36372
rect 13360 36320 13412 36372
rect 9312 36159 9364 36168
rect 9312 36125 9321 36159
rect 9321 36125 9355 36159
rect 9355 36125 9364 36159
rect 9312 36116 9364 36125
rect 756 36048 808 36100
rect 5816 36048 5868 36100
rect 6828 36048 6880 36100
rect 8300 36048 8352 36100
rect 11796 36116 11848 36168
rect 7196 35980 7248 36032
rect 12164 36116 12216 36168
rect 14188 36159 14240 36168
rect 14188 36125 14197 36159
rect 14197 36125 14231 36159
rect 14231 36125 14240 36159
rect 14188 36116 14240 36125
rect 12716 36048 12768 36100
rect 12992 36091 13044 36100
rect 12992 36057 13001 36091
rect 13001 36057 13035 36091
rect 13035 36057 13044 36091
rect 12992 36048 13044 36057
rect 13176 36048 13228 36100
rect 15568 36048 15620 36100
rect 12072 36023 12124 36032
rect 12072 35989 12081 36023
rect 12081 35989 12115 36023
rect 12115 35989 12124 36023
rect 12072 35980 12124 35989
rect 13268 36023 13320 36032
rect 13268 35989 13277 36023
rect 13277 35989 13311 36023
rect 13311 35989 13320 36023
rect 13268 35980 13320 35989
rect 15108 35980 15160 36032
rect 4376 35878 4428 35930
rect 4440 35878 4492 35930
rect 4504 35878 4556 35930
rect 4568 35878 4620 35930
rect 4632 35878 4684 35930
rect 7803 35878 7855 35930
rect 7867 35878 7919 35930
rect 7931 35878 7983 35930
rect 7995 35878 8047 35930
rect 8059 35878 8111 35930
rect 11230 35878 11282 35930
rect 11294 35878 11346 35930
rect 11358 35878 11410 35930
rect 11422 35878 11474 35930
rect 11486 35878 11538 35930
rect 14657 35878 14709 35930
rect 14721 35878 14773 35930
rect 14785 35878 14837 35930
rect 14849 35878 14901 35930
rect 14913 35878 14965 35930
rect 1768 35819 1820 35828
rect 1768 35785 1777 35819
rect 1777 35785 1811 35819
rect 1811 35785 1820 35819
rect 1768 35776 1820 35785
rect 9312 35776 9364 35828
rect 10140 35819 10192 35828
rect 10140 35785 10149 35819
rect 10149 35785 10183 35819
rect 10183 35785 10192 35819
rect 10140 35776 10192 35785
rect 10232 35708 10284 35760
rect 756 35640 808 35692
rect 1952 35683 2004 35692
rect 1952 35649 1961 35683
rect 1961 35649 1995 35683
rect 1995 35649 2004 35683
rect 1952 35640 2004 35649
rect 8576 35683 8628 35692
rect 8576 35649 8585 35683
rect 8585 35649 8619 35683
rect 8619 35649 8628 35683
rect 8576 35640 8628 35649
rect 10324 35683 10376 35692
rect 10324 35649 10333 35683
rect 10333 35649 10367 35683
rect 10367 35649 10376 35683
rect 10324 35640 10376 35649
rect 11888 35640 11940 35692
rect 12072 35640 12124 35692
rect 12440 35751 12492 35760
rect 12440 35717 12449 35751
rect 12449 35717 12483 35751
rect 12483 35717 12492 35751
rect 12440 35708 12492 35717
rect 14188 35776 14240 35828
rect 6000 35436 6052 35488
rect 13176 35572 13228 35624
rect 13544 35683 13596 35692
rect 13544 35649 13553 35683
rect 13553 35649 13587 35683
rect 13587 35649 13596 35683
rect 13544 35640 13596 35649
rect 13636 35640 13688 35692
rect 14464 35572 14516 35624
rect 15108 35504 15160 35556
rect 13820 35479 13872 35488
rect 13820 35445 13829 35479
rect 13829 35445 13863 35479
rect 13863 35445 13872 35479
rect 13820 35436 13872 35445
rect 15476 35436 15528 35488
rect 2663 35334 2715 35386
rect 2727 35334 2779 35386
rect 2791 35334 2843 35386
rect 2855 35334 2907 35386
rect 2919 35334 2971 35386
rect 6090 35334 6142 35386
rect 6154 35334 6206 35386
rect 6218 35334 6270 35386
rect 6282 35334 6334 35386
rect 6346 35334 6398 35386
rect 9517 35334 9569 35386
rect 9581 35334 9633 35386
rect 9645 35334 9697 35386
rect 9709 35334 9761 35386
rect 9773 35334 9825 35386
rect 12944 35334 12996 35386
rect 13008 35334 13060 35386
rect 13072 35334 13124 35386
rect 13136 35334 13188 35386
rect 13200 35334 13252 35386
rect 1952 35232 2004 35284
rect 10324 35232 10376 35284
rect 12808 35232 12860 35284
rect 6828 35096 6880 35148
rect 11060 35096 11112 35148
rect 11520 35139 11572 35148
rect 11520 35105 11529 35139
rect 11529 35105 11563 35139
rect 11563 35105 11572 35139
rect 11520 35096 11572 35105
rect 5540 35028 5592 35080
rect 10968 35028 11020 35080
rect 6920 34960 6972 35012
rect 11152 34960 11204 35012
rect 12164 35028 12216 35080
rect 10416 34892 10468 34944
rect 14556 34960 14608 35012
rect 12348 34892 12400 34944
rect 12532 34935 12584 34944
rect 12532 34901 12541 34935
rect 12541 34901 12575 34935
rect 12575 34901 12584 34935
rect 12532 34892 12584 34901
rect 13268 34935 13320 34944
rect 13268 34901 13277 34935
rect 13277 34901 13311 34935
rect 13311 34901 13320 34935
rect 13268 34892 13320 34901
rect 4376 34790 4428 34842
rect 4440 34790 4492 34842
rect 4504 34790 4556 34842
rect 4568 34790 4620 34842
rect 4632 34790 4684 34842
rect 7803 34790 7855 34842
rect 7867 34790 7919 34842
rect 7931 34790 7983 34842
rect 7995 34790 8047 34842
rect 8059 34790 8111 34842
rect 11230 34790 11282 34842
rect 11294 34790 11346 34842
rect 11358 34790 11410 34842
rect 11422 34790 11474 34842
rect 11486 34790 11538 34842
rect 14657 34790 14709 34842
rect 14721 34790 14773 34842
rect 14785 34790 14837 34842
rect 14849 34790 14901 34842
rect 14913 34790 14965 34842
rect 5724 34688 5776 34740
rect 6828 34688 6880 34740
rect 10416 34731 10468 34740
rect 10416 34697 10425 34731
rect 10425 34697 10459 34731
rect 10459 34697 10468 34731
rect 10416 34688 10468 34697
rect 10968 34731 11020 34740
rect 10968 34697 10977 34731
rect 10977 34697 11011 34731
rect 11011 34697 11020 34731
rect 10968 34688 11020 34697
rect 13544 34688 13596 34740
rect 11980 34620 12032 34672
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 10600 34595 10652 34604
rect 10600 34561 10609 34595
rect 10609 34561 10643 34595
rect 10643 34561 10652 34595
rect 10600 34552 10652 34561
rect 10876 34595 10928 34604
rect 10876 34561 10885 34595
rect 10885 34561 10919 34595
rect 10919 34561 10928 34595
rect 10876 34552 10928 34561
rect 11060 34552 11112 34604
rect 10508 34484 10560 34536
rect 12256 34595 12308 34604
rect 12256 34561 12265 34595
rect 12265 34561 12299 34595
rect 12299 34561 12308 34595
rect 12256 34552 12308 34561
rect 12440 34595 12492 34604
rect 12440 34561 12449 34595
rect 12449 34561 12483 34595
rect 12483 34561 12492 34595
rect 12440 34552 12492 34561
rect 13360 34595 13412 34604
rect 13360 34561 13369 34595
rect 13369 34561 13403 34595
rect 13403 34561 13412 34595
rect 13360 34552 13412 34561
rect 13544 34595 13596 34604
rect 13544 34561 13553 34595
rect 13553 34561 13587 34595
rect 13587 34561 13596 34595
rect 13544 34552 13596 34561
rect 14096 34595 14148 34604
rect 14096 34561 14105 34595
rect 14105 34561 14139 34595
rect 14139 34561 14148 34595
rect 14096 34552 14148 34561
rect 15660 34552 15712 34604
rect 12348 34484 12400 34536
rect 13820 34391 13872 34400
rect 13820 34357 13829 34391
rect 13829 34357 13863 34391
rect 13863 34357 13872 34391
rect 13820 34348 13872 34357
rect 2663 34246 2715 34298
rect 2727 34246 2779 34298
rect 2791 34246 2843 34298
rect 2855 34246 2907 34298
rect 2919 34246 2971 34298
rect 6090 34246 6142 34298
rect 6154 34246 6206 34298
rect 6218 34246 6270 34298
rect 6282 34246 6334 34298
rect 6346 34246 6398 34298
rect 9517 34246 9569 34298
rect 9581 34246 9633 34298
rect 9645 34246 9697 34298
rect 9709 34246 9761 34298
rect 9773 34246 9825 34298
rect 12944 34246 12996 34298
rect 13008 34246 13060 34298
rect 13072 34246 13124 34298
rect 13136 34246 13188 34298
rect 13200 34246 13252 34298
rect 10232 34187 10284 34196
rect 10232 34153 10241 34187
rect 10241 34153 10275 34187
rect 10275 34153 10284 34187
rect 10232 34144 10284 34153
rect 10508 34187 10560 34196
rect 10508 34153 10517 34187
rect 10517 34153 10551 34187
rect 10551 34153 10560 34187
rect 10508 34144 10560 34153
rect 11612 34008 11664 34060
rect 756 33940 808 33992
rect 8760 33940 8812 33992
rect 11520 33940 11572 33992
rect 11796 33940 11848 33992
rect 11612 33872 11664 33924
rect 12808 33940 12860 33992
rect 12992 33940 13044 33992
rect 14280 33983 14332 33992
rect 14280 33949 14289 33983
rect 14289 33949 14323 33983
rect 14323 33949 14332 33983
rect 14280 33940 14332 33949
rect 3608 33804 3660 33856
rect 9864 33804 9916 33856
rect 10324 33804 10376 33856
rect 10508 33804 10560 33856
rect 12716 33872 12768 33924
rect 12072 33804 12124 33856
rect 13268 33804 13320 33856
rect 13544 33847 13596 33856
rect 13544 33813 13553 33847
rect 13553 33813 13587 33847
rect 13587 33813 13596 33847
rect 13544 33804 13596 33813
rect 4376 33702 4428 33754
rect 4440 33702 4492 33754
rect 4504 33702 4556 33754
rect 4568 33702 4620 33754
rect 4632 33702 4684 33754
rect 7803 33702 7855 33754
rect 7867 33702 7919 33754
rect 7931 33702 7983 33754
rect 7995 33702 8047 33754
rect 8059 33702 8111 33754
rect 11230 33702 11282 33754
rect 11294 33702 11346 33754
rect 11358 33702 11410 33754
rect 11422 33702 11474 33754
rect 11486 33702 11538 33754
rect 14657 33702 14709 33754
rect 14721 33702 14773 33754
rect 14785 33702 14837 33754
rect 14849 33702 14901 33754
rect 14913 33702 14965 33754
rect 12164 33600 12216 33652
rect 10784 33532 10836 33584
rect 11796 33507 11848 33516
rect 11796 33473 11805 33507
rect 11805 33473 11839 33507
rect 11839 33473 11848 33507
rect 11796 33464 11848 33473
rect 12164 33507 12216 33516
rect 12164 33473 12171 33507
rect 12171 33473 12205 33507
rect 12205 33473 12216 33507
rect 12164 33464 12216 33473
rect 14004 33464 14056 33516
rect 15384 33464 15436 33516
rect 11612 33396 11664 33448
rect 10140 33260 10192 33312
rect 12900 33303 12952 33312
rect 12900 33269 12909 33303
rect 12909 33269 12943 33303
rect 12943 33269 12952 33303
rect 12900 33260 12952 33269
rect 12992 33260 13044 33312
rect 14004 33260 14056 33312
rect 14188 33303 14240 33312
rect 14188 33269 14197 33303
rect 14197 33269 14231 33303
rect 14231 33269 14240 33303
rect 14188 33260 14240 33269
rect 2663 33158 2715 33210
rect 2727 33158 2779 33210
rect 2791 33158 2843 33210
rect 2855 33158 2907 33210
rect 2919 33158 2971 33210
rect 6090 33158 6142 33210
rect 6154 33158 6206 33210
rect 6218 33158 6270 33210
rect 6282 33158 6334 33210
rect 6346 33158 6398 33210
rect 9517 33158 9569 33210
rect 9581 33158 9633 33210
rect 9645 33158 9697 33210
rect 9709 33158 9761 33210
rect 9773 33158 9825 33210
rect 12944 33158 12996 33210
rect 13008 33158 13060 33210
rect 13072 33158 13124 33210
rect 13136 33158 13188 33210
rect 13200 33158 13252 33210
rect 10048 33056 10100 33108
rect 10692 33056 10744 33108
rect 11796 33056 11848 33108
rect 12440 33056 12492 33108
rect 756 32852 808 32904
rect 8944 32852 8996 32904
rect 10876 32920 10928 32972
rect 8484 32784 8536 32836
rect 6460 32716 6512 32768
rect 7288 32716 7340 32768
rect 11152 32895 11204 32904
rect 11152 32861 11161 32895
rect 11161 32861 11195 32895
rect 11195 32861 11204 32895
rect 11152 32852 11204 32861
rect 13728 32988 13780 33040
rect 14280 32988 14332 33040
rect 15568 32920 15620 32972
rect 11888 32827 11940 32836
rect 11888 32793 11897 32827
rect 11897 32793 11931 32827
rect 11931 32793 11940 32827
rect 11888 32784 11940 32793
rect 11060 32716 11112 32768
rect 11980 32716 12032 32768
rect 12164 32759 12216 32768
rect 12164 32725 12173 32759
rect 12173 32725 12207 32759
rect 12207 32725 12216 32759
rect 12164 32716 12216 32725
rect 14280 32895 14332 32904
rect 14280 32861 14289 32895
rect 14289 32861 14323 32895
rect 14323 32861 14332 32895
rect 14280 32852 14332 32861
rect 12440 32827 12492 32836
rect 12440 32793 12449 32827
rect 12449 32793 12483 32827
rect 12483 32793 12492 32827
rect 12440 32784 12492 32793
rect 12716 32784 12768 32836
rect 13360 32827 13412 32836
rect 13360 32793 13369 32827
rect 13369 32793 13403 32827
rect 13403 32793 13412 32827
rect 13360 32784 13412 32793
rect 12992 32716 13044 32768
rect 14556 32784 14608 32836
rect 4376 32614 4428 32666
rect 4440 32614 4492 32666
rect 4504 32614 4556 32666
rect 4568 32614 4620 32666
rect 4632 32614 4684 32666
rect 7803 32614 7855 32666
rect 7867 32614 7919 32666
rect 7931 32614 7983 32666
rect 7995 32614 8047 32666
rect 8059 32614 8111 32666
rect 11230 32614 11282 32666
rect 11294 32614 11346 32666
rect 11358 32614 11410 32666
rect 11422 32614 11474 32666
rect 11486 32614 11538 32666
rect 14657 32614 14709 32666
rect 14721 32614 14773 32666
rect 14785 32614 14837 32666
rect 14849 32614 14901 32666
rect 14913 32614 14965 32666
rect 2228 32512 2280 32564
rect 756 32376 808 32428
rect 2228 32419 2280 32428
rect 2228 32385 2237 32419
rect 2237 32385 2271 32419
rect 2271 32385 2280 32419
rect 2228 32376 2280 32385
rect 6920 32376 6972 32428
rect 7288 32415 7313 32428
rect 7313 32415 7340 32428
rect 7288 32376 7340 32415
rect 8668 32512 8720 32564
rect 8484 32444 8536 32496
rect 9864 32512 9916 32564
rect 12992 32512 13044 32564
rect 13544 32512 13596 32564
rect 11980 32444 12032 32496
rect 10324 32419 10376 32428
rect 10324 32385 10333 32419
rect 10333 32385 10376 32419
rect 1860 32172 1912 32224
rect 8024 32215 8076 32224
rect 8024 32181 8033 32215
rect 8033 32181 8067 32215
rect 8067 32181 8076 32215
rect 8024 32172 8076 32181
rect 10324 32376 10376 32385
rect 11060 32376 11112 32428
rect 12992 32419 13044 32428
rect 12992 32385 13001 32419
rect 13001 32385 13035 32419
rect 13035 32385 13044 32419
rect 12992 32376 13044 32385
rect 11520 32351 11572 32360
rect 9404 32215 9456 32224
rect 9404 32181 9413 32215
rect 9413 32181 9447 32215
rect 9447 32181 9456 32215
rect 9404 32172 9456 32181
rect 11520 32317 11529 32351
rect 11529 32317 11563 32351
rect 11563 32317 11572 32351
rect 11520 32308 11572 32317
rect 14096 32419 14148 32428
rect 14096 32385 14105 32419
rect 14105 32385 14139 32419
rect 14139 32385 14148 32419
rect 14096 32376 14148 32385
rect 14188 32308 14240 32360
rect 12532 32215 12584 32224
rect 12532 32181 12541 32215
rect 12541 32181 12575 32215
rect 12575 32181 12584 32215
rect 12532 32172 12584 32181
rect 12624 32172 12676 32224
rect 13544 32172 13596 32224
rect 14004 32172 14056 32224
rect 15108 32172 15160 32224
rect 2663 32070 2715 32122
rect 2727 32070 2779 32122
rect 2791 32070 2843 32122
rect 2855 32070 2907 32122
rect 2919 32070 2971 32122
rect 6090 32070 6142 32122
rect 6154 32070 6206 32122
rect 6218 32070 6270 32122
rect 6282 32070 6334 32122
rect 6346 32070 6398 32122
rect 9517 32070 9569 32122
rect 9581 32070 9633 32122
rect 9645 32070 9697 32122
rect 9709 32070 9761 32122
rect 9773 32070 9825 32122
rect 12944 32070 12996 32122
rect 13008 32070 13060 32122
rect 13072 32070 13124 32122
rect 13136 32070 13188 32122
rect 13200 32070 13252 32122
rect 6460 31968 6512 32020
rect 8300 31968 8352 32020
rect 8944 32011 8996 32020
rect 8944 31977 8953 32011
rect 8953 31977 8987 32011
rect 8987 31977 8996 32011
rect 8944 31968 8996 31977
rect 10416 31968 10468 32020
rect 10784 32011 10836 32020
rect 10784 31977 10793 32011
rect 10793 31977 10827 32011
rect 10827 31977 10836 32011
rect 10784 31968 10836 31977
rect 12348 31968 12400 32020
rect 14280 31968 14332 32020
rect 1860 31764 1912 31816
rect 6644 31832 6696 31884
rect 7196 31832 7248 31884
rect 7472 31764 7524 31816
rect 11980 31900 12032 31952
rect 12532 31900 12584 31952
rect 14004 31900 14056 31952
rect 14464 31900 14516 31952
rect 13820 31875 13872 31884
rect 13820 31841 13829 31875
rect 13829 31841 13863 31875
rect 13863 31841 13872 31875
rect 13820 31832 13872 31841
rect 10784 31764 10836 31816
rect 6920 31696 6972 31748
rect 7196 31696 7248 31748
rect 10876 31696 10928 31748
rect 11520 31807 11572 31816
rect 11520 31773 11529 31807
rect 11529 31773 11563 31807
rect 11563 31773 11572 31807
rect 11520 31764 11572 31773
rect 11612 31764 11664 31816
rect 11980 31807 12032 31816
rect 11980 31773 11989 31807
rect 11989 31773 12023 31807
rect 12023 31773 12032 31807
rect 11980 31764 12032 31773
rect 12348 31764 12400 31816
rect 12900 31807 12952 31816
rect 12900 31773 12909 31807
rect 12909 31773 12943 31807
rect 12943 31773 12952 31807
rect 12900 31764 12952 31773
rect 13084 31764 13136 31816
rect 13176 31807 13228 31816
rect 13176 31773 13185 31807
rect 13185 31773 13219 31807
rect 13219 31773 13228 31807
rect 13176 31764 13228 31773
rect 14280 31807 14332 31816
rect 14280 31773 14289 31807
rect 14289 31773 14323 31807
rect 14323 31773 14332 31807
rect 14280 31764 14332 31773
rect 6552 31628 6604 31680
rect 9128 31628 9180 31680
rect 9312 31628 9364 31680
rect 13452 31628 13504 31680
rect 4376 31526 4428 31578
rect 4440 31526 4492 31578
rect 4504 31526 4556 31578
rect 4568 31526 4620 31578
rect 4632 31526 4684 31578
rect 7803 31526 7855 31578
rect 7867 31526 7919 31578
rect 7931 31526 7983 31578
rect 7995 31526 8047 31578
rect 8059 31526 8111 31578
rect 11230 31526 11282 31578
rect 11294 31526 11346 31578
rect 11358 31526 11410 31578
rect 11422 31526 11474 31578
rect 11486 31526 11538 31578
rect 14657 31526 14709 31578
rect 14721 31526 14773 31578
rect 14785 31526 14837 31578
rect 14849 31526 14901 31578
rect 14913 31526 14965 31578
rect 10784 31424 10836 31476
rect 10876 31424 10928 31476
rect 11888 31424 11940 31476
rect 6644 31356 6696 31408
rect 7564 31356 7616 31408
rect 9036 31356 9088 31408
rect 756 31288 808 31340
rect 2228 31288 2280 31340
rect 6828 31288 6880 31340
rect 8484 31288 8536 31340
rect 10140 31288 10192 31340
rect 10876 31331 10928 31340
rect 10876 31297 10885 31331
rect 10885 31297 10919 31331
rect 10919 31297 10928 31331
rect 10876 31288 10928 31297
rect 13452 31356 13504 31408
rect 11888 31288 11940 31340
rect 12716 31331 12768 31340
rect 12716 31297 12725 31331
rect 12725 31297 12759 31331
rect 12759 31297 12768 31331
rect 12716 31288 12768 31297
rect 14096 31331 14148 31340
rect 14096 31297 14105 31331
rect 14105 31297 14139 31331
rect 14139 31297 14148 31331
rect 14096 31288 14148 31297
rect 11244 31220 11296 31272
rect 12164 31263 12216 31272
rect 12164 31229 12173 31263
rect 12173 31229 12207 31263
rect 12207 31229 12216 31263
rect 12164 31220 12216 31229
rect 12440 31263 12492 31272
rect 12440 31229 12449 31263
rect 12449 31229 12483 31263
rect 12483 31229 12492 31263
rect 12440 31220 12492 31229
rect 12532 31263 12584 31272
rect 12532 31229 12566 31263
rect 12566 31229 12584 31263
rect 12532 31220 12584 31229
rect 13268 31220 13320 31272
rect 13636 31220 13688 31272
rect 11888 31152 11940 31204
rect 1216 31084 1268 31136
rect 10416 31084 10468 31136
rect 10784 31084 10836 31136
rect 12532 31084 12584 31136
rect 13820 31127 13872 31136
rect 13820 31093 13829 31127
rect 13829 31093 13863 31127
rect 13863 31093 13872 31127
rect 13820 31084 13872 31093
rect 15752 31084 15804 31136
rect 2663 30982 2715 31034
rect 2727 30982 2779 31034
rect 2791 30982 2843 31034
rect 2855 30982 2907 31034
rect 2919 30982 2971 31034
rect 6090 30982 6142 31034
rect 6154 30982 6206 31034
rect 6218 30982 6270 31034
rect 6282 30982 6334 31034
rect 6346 30982 6398 31034
rect 9517 30982 9569 31034
rect 9581 30982 9633 31034
rect 9645 30982 9697 31034
rect 9709 30982 9761 31034
rect 9773 30982 9825 31034
rect 12944 30982 12996 31034
rect 13008 30982 13060 31034
rect 13072 30982 13124 31034
rect 13136 30982 13188 31034
rect 13200 30982 13252 31034
rect 6736 30880 6788 30932
rect 10876 30880 10928 30932
rect 13912 30923 13964 30932
rect 13912 30889 13921 30923
rect 13921 30889 13955 30923
rect 13955 30889 13964 30923
rect 13912 30880 13964 30889
rect 10324 30812 10376 30864
rect 7012 30744 7064 30796
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 8668 30744 8720 30796
rect 8852 30744 8904 30796
rect 11796 30744 11848 30796
rect 10508 30676 10560 30728
rect 12716 30855 12768 30864
rect 12716 30821 12725 30855
rect 12725 30821 12759 30855
rect 12759 30821 12768 30855
rect 12716 30812 12768 30821
rect 12624 30744 12676 30796
rect 12808 30744 12860 30796
rect 13636 30744 13688 30796
rect 11060 30651 11112 30660
rect 11060 30617 11069 30651
rect 11069 30617 11103 30651
rect 11103 30617 11112 30651
rect 11060 30608 11112 30617
rect 11980 30651 12032 30660
rect 11980 30617 11989 30651
rect 11989 30617 12023 30651
rect 12023 30617 12032 30651
rect 11980 30608 12032 30617
rect 13176 30676 13228 30728
rect 5264 30540 5316 30592
rect 7288 30540 7340 30592
rect 8392 30540 8444 30592
rect 8668 30540 8720 30592
rect 10140 30540 10192 30592
rect 12072 30540 12124 30592
rect 12440 30540 12492 30592
rect 4376 30438 4428 30490
rect 4440 30438 4492 30490
rect 4504 30438 4556 30490
rect 4568 30438 4620 30490
rect 4632 30438 4684 30490
rect 7803 30438 7855 30490
rect 7867 30438 7919 30490
rect 7931 30438 7983 30490
rect 7995 30438 8047 30490
rect 8059 30438 8111 30490
rect 11230 30438 11282 30490
rect 11294 30438 11346 30490
rect 11358 30438 11410 30490
rect 11422 30438 11474 30490
rect 11486 30438 11538 30490
rect 14657 30438 14709 30490
rect 14721 30438 14773 30490
rect 14785 30438 14837 30490
rect 14849 30438 14901 30490
rect 14913 30438 14965 30490
rect 6644 30336 6696 30388
rect 8576 30336 8628 30388
rect 9312 30336 9364 30388
rect 9496 30336 9548 30388
rect 10876 30336 10928 30388
rect 7472 30268 7524 30320
rect 6552 30200 6604 30252
rect 7012 30200 7064 30252
rect 9404 30243 9456 30252
rect 9404 30209 9413 30243
rect 9413 30209 9447 30243
rect 9447 30209 9456 30243
rect 9404 30200 9456 30209
rect 10876 30200 10928 30252
rect 11336 30311 11388 30320
rect 11336 30277 11345 30311
rect 11345 30277 11379 30311
rect 11379 30277 11388 30311
rect 11336 30268 11388 30277
rect 11520 30200 11572 30252
rect 8116 30132 8168 30184
rect 8484 30132 8536 30184
rect 9312 30132 9364 30184
rect 10140 30132 10192 30184
rect 12256 30200 12308 30252
rect 8944 30064 8996 30116
rect 11152 30064 11204 30116
rect 7288 29996 7340 30048
rect 9956 29996 10008 30048
rect 10968 29996 11020 30048
rect 11244 29996 11296 30048
rect 15568 30200 15620 30252
rect 15476 30132 15528 30184
rect 13912 30064 13964 30116
rect 12164 29996 12216 30048
rect 12624 29996 12676 30048
rect 12900 30039 12952 30048
rect 12900 30005 12909 30039
rect 12909 30005 12943 30039
rect 12943 30005 12952 30039
rect 12900 29996 12952 30005
rect 14556 29996 14608 30048
rect 15108 29996 15160 30048
rect 15568 29996 15620 30048
rect 2663 29894 2715 29946
rect 2727 29894 2779 29946
rect 2791 29894 2843 29946
rect 2855 29894 2907 29946
rect 2919 29894 2971 29946
rect 6090 29894 6142 29946
rect 6154 29894 6206 29946
rect 6218 29894 6270 29946
rect 6282 29894 6334 29946
rect 6346 29894 6398 29946
rect 9517 29894 9569 29946
rect 9581 29894 9633 29946
rect 9645 29894 9697 29946
rect 9709 29894 9761 29946
rect 9773 29894 9825 29946
rect 12944 29894 12996 29946
rect 13008 29894 13060 29946
rect 13072 29894 13124 29946
rect 13136 29894 13188 29946
rect 13200 29894 13252 29946
rect 8116 29792 8168 29844
rect 10048 29792 10100 29844
rect 9956 29724 10008 29776
rect 10692 29792 10744 29844
rect 10784 29792 10836 29844
rect 8576 29656 8628 29708
rect 756 29588 808 29640
rect 10140 29588 10192 29640
rect 11336 29767 11388 29776
rect 11336 29733 11345 29767
rect 11345 29733 11379 29767
rect 11379 29733 11388 29767
rect 11336 29724 11388 29733
rect 12624 29792 12676 29844
rect 13544 29724 13596 29776
rect 11244 29588 11296 29640
rect 11428 29588 11480 29640
rect 12624 29656 12676 29708
rect 13728 29588 13780 29640
rect 8576 29520 8628 29572
rect 1768 29452 1820 29504
rect 8760 29452 8812 29504
rect 9956 29495 10008 29504
rect 9956 29461 9965 29495
rect 9965 29461 9999 29495
rect 9999 29461 10008 29495
rect 9956 29452 10008 29461
rect 11336 29520 11388 29572
rect 12992 29520 13044 29572
rect 13544 29563 13596 29572
rect 13544 29529 13553 29563
rect 13553 29529 13587 29563
rect 13587 29529 13596 29563
rect 13544 29520 13596 29529
rect 12624 29452 12676 29504
rect 13636 29495 13688 29504
rect 13636 29461 13645 29495
rect 13645 29461 13679 29495
rect 13679 29461 13688 29495
rect 13636 29452 13688 29461
rect 4376 29350 4428 29402
rect 4440 29350 4492 29402
rect 4504 29350 4556 29402
rect 4568 29350 4620 29402
rect 4632 29350 4684 29402
rect 7803 29350 7855 29402
rect 7867 29350 7919 29402
rect 7931 29350 7983 29402
rect 7995 29350 8047 29402
rect 8059 29350 8111 29402
rect 11230 29350 11282 29402
rect 11294 29350 11346 29402
rect 11358 29350 11410 29402
rect 11422 29350 11474 29402
rect 11486 29350 11538 29402
rect 14657 29350 14709 29402
rect 14721 29350 14773 29402
rect 14785 29350 14837 29402
rect 14849 29350 14901 29402
rect 14913 29350 14965 29402
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 2412 29112 2464 29164
rect 8484 29248 8536 29300
rect 8760 29248 8812 29300
rect 9864 29291 9916 29300
rect 9864 29257 9873 29291
rect 9873 29257 9907 29291
rect 9907 29257 9916 29291
rect 9864 29248 9916 29257
rect 11244 29248 11296 29300
rect 11060 29180 11112 29232
rect 9220 29155 9272 29164
rect 9220 29121 9229 29155
rect 9229 29121 9263 29155
rect 9263 29121 9272 29155
rect 9220 29112 9272 29121
rect 12256 29248 12308 29300
rect 12624 29248 12676 29300
rect 7012 29044 7064 29096
rect 8392 29044 8444 29096
rect 8944 29087 8996 29096
rect 1952 28976 2004 29028
rect 7288 28976 7340 29028
rect 8944 29053 8953 29087
rect 8953 29053 8987 29087
rect 8987 29053 8996 29087
rect 8944 29044 8996 29053
rect 8208 28908 8260 28960
rect 9864 29044 9916 29096
rect 12162 29155 12214 29164
rect 12162 29121 12173 29155
rect 12173 29121 12207 29155
rect 12207 29121 12214 29155
rect 12162 29112 12214 29121
rect 11244 28976 11296 29028
rect 11520 28976 11572 29028
rect 11060 28951 11112 28960
rect 11060 28917 11069 28951
rect 11069 28917 11103 28951
rect 11103 28917 11112 28951
rect 11060 28908 11112 28917
rect 12256 28908 12308 28960
rect 12992 29044 13044 29096
rect 13176 29087 13228 29096
rect 13176 29053 13185 29087
rect 13185 29053 13219 29087
rect 13219 29053 13228 29087
rect 13176 29044 13228 29053
rect 14188 29112 14240 29164
rect 15108 28976 15160 29028
rect 12716 28908 12768 28960
rect 13544 28908 13596 28960
rect 2663 28806 2715 28858
rect 2727 28806 2779 28858
rect 2791 28806 2843 28858
rect 2855 28806 2907 28858
rect 2919 28806 2971 28858
rect 6090 28806 6142 28858
rect 6154 28806 6206 28858
rect 6218 28806 6270 28858
rect 6282 28806 6334 28858
rect 6346 28806 6398 28858
rect 9517 28806 9569 28858
rect 9581 28806 9633 28858
rect 9645 28806 9697 28858
rect 9709 28806 9761 28858
rect 9773 28806 9825 28858
rect 12944 28806 12996 28858
rect 13008 28806 13060 28858
rect 13072 28806 13124 28858
rect 13136 28806 13188 28858
rect 13200 28806 13252 28858
rect 6828 28704 6880 28756
rect 7380 28704 7432 28756
rect 8760 28704 8812 28756
rect 9312 28636 9364 28688
rect 1216 28500 1268 28552
rect 6644 28543 6696 28552
rect 6644 28509 6651 28543
rect 6651 28509 6685 28543
rect 6685 28509 6696 28543
rect 6644 28500 6696 28509
rect 9036 28500 9088 28552
rect 9588 28704 9640 28756
rect 10324 28704 10376 28756
rect 13728 28704 13780 28756
rect 14004 28704 14056 28756
rect 9956 28636 10008 28688
rect 9496 28568 9548 28620
rect 10416 28611 10468 28620
rect 10416 28577 10425 28611
rect 10425 28577 10459 28611
rect 10459 28577 10468 28611
rect 10416 28568 10468 28577
rect 12624 28636 12676 28688
rect 12808 28636 12860 28688
rect 13176 28568 13228 28620
rect 13820 28568 13872 28620
rect 9588 28500 9640 28552
rect 10324 28500 10376 28552
rect 12072 28543 12124 28552
rect 12072 28509 12081 28543
rect 12081 28509 12115 28543
rect 12115 28509 12124 28543
rect 12072 28500 12124 28509
rect 12992 28543 13044 28552
rect 12992 28509 13001 28543
rect 13001 28509 13035 28543
rect 13035 28509 13044 28543
rect 12992 28500 13044 28509
rect 7472 28364 7524 28416
rect 10692 28364 10744 28416
rect 11520 28364 11572 28416
rect 11888 28407 11940 28416
rect 11888 28373 11897 28407
rect 11897 28373 11931 28407
rect 11931 28373 11940 28407
rect 11888 28364 11940 28373
rect 13360 28364 13412 28416
rect 4376 28262 4428 28314
rect 4440 28262 4492 28314
rect 4504 28262 4556 28314
rect 4568 28262 4620 28314
rect 4632 28262 4684 28314
rect 7803 28262 7855 28314
rect 7867 28262 7919 28314
rect 7931 28262 7983 28314
rect 7995 28262 8047 28314
rect 8059 28262 8111 28314
rect 11230 28262 11282 28314
rect 11294 28262 11346 28314
rect 11358 28262 11410 28314
rect 11422 28262 11474 28314
rect 11486 28262 11538 28314
rect 14657 28262 14709 28314
rect 14721 28262 14773 28314
rect 14785 28262 14837 28314
rect 14849 28262 14901 28314
rect 14913 28262 14965 28314
rect 1400 28160 1452 28212
rect 7380 28160 7432 28212
rect 7564 28097 7616 28144
rect 756 28024 808 28076
rect 6828 28024 6880 28076
rect 7564 28092 7589 28097
rect 7589 28092 7616 28097
rect 9588 28160 9640 28212
rect 9956 28160 10008 28212
rect 10324 28160 10376 28212
rect 10508 28203 10560 28212
rect 10508 28169 10517 28203
rect 10517 28169 10551 28203
rect 10551 28169 10560 28203
rect 10508 28160 10560 28169
rect 12256 28160 12308 28212
rect 7104 27820 7156 27872
rect 9772 28024 9824 28076
rect 9036 27956 9088 28008
rect 9404 27956 9456 28008
rect 9864 27999 9916 28008
rect 9864 27965 9873 27999
rect 9873 27965 9907 27999
rect 9907 27965 9916 27999
rect 9864 27956 9916 27965
rect 8116 27820 8168 27872
rect 8484 27820 8536 27872
rect 11060 27888 11112 27940
rect 12716 28024 12768 28076
rect 13820 28092 13872 28144
rect 13544 28024 13596 28076
rect 15568 28024 15620 28076
rect 11520 27956 11572 28008
rect 11612 27888 11664 27940
rect 12532 27820 12584 27872
rect 12808 27863 12860 27872
rect 12808 27829 12817 27863
rect 12817 27829 12851 27863
rect 12851 27829 12860 27863
rect 12808 27820 12860 27829
rect 13176 27820 13228 27872
rect 13544 27820 13596 27872
rect 13912 27820 13964 27872
rect 2663 27718 2715 27770
rect 2727 27718 2779 27770
rect 2791 27718 2843 27770
rect 2855 27718 2907 27770
rect 2919 27718 2971 27770
rect 6090 27718 6142 27770
rect 6154 27718 6206 27770
rect 6218 27718 6270 27770
rect 6282 27718 6334 27770
rect 6346 27718 6398 27770
rect 9517 27718 9569 27770
rect 9581 27718 9633 27770
rect 9645 27718 9697 27770
rect 9709 27718 9761 27770
rect 9773 27718 9825 27770
rect 12944 27718 12996 27770
rect 13008 27718 13060 27770
rect 13072 27718 13124 27770
rect 13136 27718 13188 27770
rect 13200 27718 13252 27770
rect 6828 27480 6880 27532
rect 7288 27616 7340 27668
rect 9864 27616 9916 27668
rect 12072 27616 12124 27668
rect 15844 27616 15896 27668
rect 11612 27548 11664 27600
rect 13452 27548 13504 27600
rect 13636 27548 13688 27600
rect 7840 27480 7892 27532
rect 8116 27480 8168 27532
rect 8944 27523 8996 27532
rect 8944 27489 8953 27523
rect 8953 27489 8987 27523
rect 8987 27489 8996 27523
rect 8944 27480 8996 27489
rect 10140 27480 10192 27532
rect 10324 27480 10376 27532
rect 11704 27480 11756 27532
rect 4896 27455 4948 27464
rect 4896 27421 4905 27455
rect 4905 27421 4939 27455
rect 4939 27421 4948 27455
rect 4896 27412 4948 27421
rect 756 27344 808 27396
rect 5264 27344 5316 27396
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 9220 27455 9272 27464
rect 9220 27421 9229 27455
rect 9229 27421 9272 27455
rect 9220 27412 9272 27421
rect 12164 27480 12216 27532
rect 12440 27480 12492 27532
rect 13452 27412 13504 27464
rect 10140 27344 10192 27396
rect 6736 27276 6788 27328
rect 6828 27276 6880 27328
rect 8208 27276 8260 27328
rect 11152 27319 11204 27328
rect 11152 27285 11161 27319
rect 11161 27285 11195 27319
rect 11195 27285 11204 27319
rect 11152 27276 11204 27285
rect 11704 27319 11756 27328
rect 11704 27285 11713 27319
rect 11713 27285 11747 27319
rect 11747 27285 11756 27319
rect 11704 27276 11756 27285
rect 14188 27344 14240 27396
rect 13268 27276 13320 27328
rect 13820 27276 13872 27328
rect 4376 27174 4428 27226
rect 4440 27174 4492 27226
rect 4504 27174 4556 27226
rect 4568 27174 4620 27226
rect 4632 27174 4684 27226
rect 7803 27174 7855 27226
rect 7867 27174 7919 27226
rect 7931 27174 7983 27226
rect 7995 27174 8047 27226
rect 8059 27174 8111 27226
rect 11230 27174 11282 27226
rect 11294 27174 11346 27226
rect 11358 27174 11410 27226
rect 11422 27174 11474 27226
rect 11486 27174 11538 27226
rect 14657 27174 14709 27226
rect 14721 27174 14773 27226
rect 14785 27174 14837 27226
rect 14849 27174 14901 27226
rect 14913 27174 14965 27226
rect 3056 27072 3108 27124
rect 3056 26936 3108 26988
rect 4160 26936 4212 26988
rect 8576 27115 8628 27124
rect 8576 27081 8585 27115
rect 8585 27081 8619 27115
rect 8619 27081 8628 27115
rect 8576 27072 8628 27081
rect 8852 27072 8904 27124
rect 11704 27072 11756 27124
rect 14648 27072 14700 27124
rect 10692 27004 10744 27056
rect 10968 27004 11020 27056
rect 5908 26936 5960 26988
rect 6460 26936 6512 26988
rect 8576 26936 8628 26988
rect 11428 26936 11480 26988
rect 13360 27047 13412 27056
rect 13360 27013 13369 27047
rect 13369 27013 13403 27047
rect 13403 27013 13412 27047
rect 13360 27004 13412 27013
rect 13728 27047 13780 27056
rect 13728 27013 13737 27047
rect 13737 27013 13771 27047
rect 13771 27013 13780 27047
rect 13728 27004 13780 27013
rect 14096 27004 14148 27056
rect 12440 26979 12492 26988
rect 12440 26945 12449 26979
rect 12449 26945 12483 26979
rect 12483 26945 12492 26979
rect 12440 26936 12492 26945
rect 12716 26979 12768 26988
rect 12716 26945 12725 26979
rect 12725 26945 12759 26979
rect 12759 26945 12768 26979
rect 12716 26936 12768 26945
rect 4896 26911 4948 26920
rect 4896 26877 4905 26911
rect 4905 26877 4939 26911
rect 4939 26877 4948 26911
rect 4896 26868 4948 26877
rect 6736 26911 6788 26920
rect 6736 26877 6745 26911
rect 6745 26877 6779 26911
rect 6779 26877 6788 26911
rect 6736 26868 6788 26877
rect 6828 26868 6880 26920
rect 7104 26732 7156 26784
rect 7748 26911 7800 26920
rect 7748 26877 7782 26911
rect 7782 26877 7800 26911
rect 7748 26868 7800 26877
rect 7932 26911 7984 26920
rect 7932 26877 7941 26911
rect 7941 26877 7975 26911
rect 7975 26877 7984 26911
rect 7932 26868 7984 26877
rect 8944 26868 8996 26920
rect 9864 26868 9916 26920
rect 11704 26911 11756 26920
rect 11704 26877 11713 26911
rect 11713 26877 11747 26911
rect 11747 26877 11756 26911
rect 11704 26868 11756 26877
rect 9036 26800 9088 26852
rect 13176 26800 13228 26852
rect 13360 26800 13412 26852
rect 11520 26732 11572 26784
rect 12716 26732 12768 26784
rect 14004 26775 14056 26784
rect 14004 26741 14013 26775
rect 14013 26741 14047 26775
rect 14047 26741 14056 26775
rect 14004 26732 14056 26741
rect 14096 26732 14148 26784
rect 2663 26630 2715 26682
rect 2727 26630 2779 26682
rect 2791 26630 2843 26682
rect 2855 26630 2907 26682
rect 2919 26630 2971 26682
rect 6090 26630 6142 26682
rect 6154 26630 6206 26682
rect 6218 26630 6270 26682
rect 6282 26630 6334 26682
rect 6346 26630 6398 26682
rect 9517 26630 9569 26682
rect 9581 26630 9633 26682
rect 9645 26630 9697 26682
rect 9709 26630 9761 26682
rect 9773 26630 9825 26682
rect 12944 26630 12996 26682
rect 13008 26630 13060 26682
rect 13072 26630 13124 26682
rect 13136 26630 13188 26682
rect 13200 26630 13252 26682
rect 3056 26528 3108 26580
rect 3056 26367 3108 26376
rect 3056 26333 3065 26367
rect 3065 26333 3099 26367
rect 3099 26333 3108 26367
rect 3056 26324 3108 26333
rect 7104 26528 7156 26580
rect 7932 26528 7984 26580
rect 10968 26528 11020 26580
rect 11428 26528 11480 26580
rect 11520 26571 11572 26580
rect 11520 26537 11529 26571
rect 11529 26537 11563 26571
rect 11563 26537 11572 26571
rect 11520 26528 11572 26537
rect 13268 26528 13320 26580
rect 12072 26460 12124 26512
rect 12440 26460 12492 26512
rect 12808 26460 12860 26512
rect 7472 26392 7524 26444
rect 9864 26392 9916 26444
rect 10232 26324 10284 26376
rect 12624 26392 12676 26444
rect 13912 26392 13964 26444
rect 1492 26299 1544 26308
rect 1492 26265 1501 26299
rect 1501 26265 1535 26299
rect 1535 26265 1544 26299
rect 1492 26256 1544 26265
rect 1584 26256 1636 26308
rect 8576 26256 8628 26308
rect 8760 26256 8812 26308
rect 12164 26324 12216 26376
rect 12440 26324 12492 26376
rect 13176 26324 13228 26376
rect 15476 26188 15528 26240
rect 15752 26188 15804 26240
rect 4376 26086 4428 26138
rect 4440 26086 4492 26138
rect 4504 26086 4556 26138
rect 4568 26086 4620 26138
rect 4632 26086 4684 26138
rect 7803 26086 7855 26138
rect 7867 26086 7919 26138
rect 7931 26086 7983 26138
rect 7995 26086 8047 26138
rect 8059 26086 8111 26138
rect 11230 26086 11282 26138
rect 11294 26086 11346 26138
rect 11358 26086 11410 26138
rect 11422 26086 11474 26138
rect 11486 26086 11538 26138
rect 14657 26086 14709 26138
rect 14721 26086 14773 26138
rect 14785 26086 14837 26138
rect 14849 26086 14901 26138
rect 14913 26086 14965 26138
rect 5080 25916 5132 25968
rect 13360 25984 13412 26036
rect 14096 25984 14148 26036
rect 4160 25848 4212 25900
rect 10232 25848 10284 25900
rect 12992 25848 13044 25900
rect 13820 25891 13872 25900
rect 13820 25857 13829 25891
rect 13829 25857 13863 25891
rect 13863 25857 13872 25891
rect 13820 25848 13872 25857
rect 756 25780 808 25832
rect 9220 25780 9272 25832
rect 10692 25780 10744 25832
rect 10968 25780 11020 25832
rect 12164 25780 12216 25832
rect 12440 25780 12492 25832
rect 13176 25780 13228 25832
rect 13544 25823 13596 25832
rect 13544 25789 13553 25823
rect 13553 25789 13587 25823
rect 13587 25789 13596 25823
rect 13544 25780 13596 25789
rect 13636 25780 13688 25832
rect 12808 25712 12860 25764
rect 13268 25755 13320 25764
rect 13268 25721 13277 25755
rect 13277 25721 13311 25755
rect 13311 25721 13320 25755
rect 13268 25712 13320 25721
rect 10968 25644 11020 25696
rect 11888 25687 11940 25696
rect 11888 25653 11897 25687
rect 11897 25653 11931 25687
rect 11931 25653 11940 25687
rect 11888 25644 11940 25653
rect 14188 25644 14240 25696
rect 2663 25542 2715 25594
rect 2727 25542 2779 25594
rect 2791 25542 2843 25594
rect 2855 25542 2907 25594
rect 2919 25542 2971 25594
rect 6090 25542 6142 25594
rect 6154 25542 6206 25594
rect 6218 25542 6270 25594
rect 6282 25542 6334 25594
rect 6346 25542 6398 25594
rect 9517 25542 9569 25594
rect 9581 25542 9633 25594
rect 9645 25542 9697 25594
rect 9709 25542 9761 25594
rect 9773 25542 9825 25594
rect 12944 25542 12996 25594
rect 13008 25542 13060 25594
rect 13072 25542 13124 25594
rect 13136 25542 13188 25594
rect 13200 25542 13252 25594
rect 10600 25440 10652 25492
rect 10784 25483 10836 25492
rect 10784 25449 10793 25483
rect 10793 25449 10827 25483
rect 10827 25449 10836 25483
rect 10784 25440 10836 25449
rect 9496 25304 9548 25356
rect 12348 25440 12400 25492
rect 13268 25440 13320 25492
rect 14556 25372 14608 25424
rect 15568 25372 15620 25424
rect 7104 25236 7156 25288
rect 7380 25236 7432 25288
rect 8208 25236 8260 25288
rect 8484 25236 8536 25288
rect 9864 25279 9916 25288
rect 9864 25245 9873 25279
rect 9873 25245 9907 25279
rect 9907 25245 9916 25279
rect 9864 25236 9916 25245
rect 9956 25279 10008 25288
rect 9956 25245 9990 25279
rect 9990 25245 10008 25279
rect 9956 25236 10008 25245
rect 8208 25100 8260 25152
rect 11980 25168 12032 25220
rect 13544 25211 13596 25220
rect 13544 25177 13553 25211
rect 13553 25177 13587 25211
rect 13587 25177 13596 25211
rect 13544 25168 13596 25177
rect 13912 25211 13964 25220
rect 13912 25177 13921 25211
rect 13921 25177 13955 25211
rect 13955 25177 13964 25211
rect 13912 25168 13964 25177
rect 4376 24998 4428 25050
rect 4440 24998 4492 25050
rect 4504 24998 4556 25050
rect 4568 24998 4620 25050
rect 4632 24998 4684 25050
rect 7803 24998 7855 25050
rect 7867 24998 7919 25050
rect 7931 24998 7983 25050
rect 7995 24998 8047 25050
rect 8059 24998 8111 25050
rect 11230 24998 11282 25050
rect 11294 24998 11346 25050
rect 11358 24998 11410 25050
rect 11422 24998 11474 25050
rect 11486 24998 11538 25050
rect 14657 24998 14709 25050
rect 14721 24998 14773 25050
rect 14785 24998 14837 25050
rect 14849 24998 14901 25050
rect 14913 24998 14965 25050
rect 7196 24896 7248 24948
rect 7748 24896 7800 24948
rect 9496 24939 9548 24948
rect 9496 24905 9505 24939
rect 9505 24905 9539 24939
rect 9539 24905 9548 24939
rect 9496 24896 9548 24905
rect 9864 24896 9916 24948
rect 11244 24896 11296 24948
rect 12072 24896 12124 24948
rect 6552 24828 6604 24880
rect 756 24760 808 24812
rect 5908 24692 5960 24744
rect 6644 24760 6696 24812
rect 7380 24760 7432 24812
rect 7564 24760 7616 24812
rect 8760 24803 8812 24812
rect 8760 24769 8769 24803
rect 8769 24769 8812 24803
rect 8760 24760 8812 24769
rect 10416 24760 10468 24812
rect 13176 24803 13228 24812
rect 13176 24769 13183 24803
rect 13183 24769 13217 24803
rect 13217 24769 13228 24803
rect 13176 24760 13228 24769
rect 7932 24692 7984 24744
rect 9220 24692 9272 24744
rect 5540 24624 5592 24676
rect 7380 24624 7432 24676
rect 8392 24624 8444 24676
rect 7472 24599 7524 24608
rect 7472 24565 7481 24599
rect 7481 24565 7515 24599
rect 7515 24565 7524 24599
rect 7472 24556 7524 24565
rect 7840 24556 7892 24608
rect 8944 24556 8996 24608
rect 9864 24556 9916 24608
rect 11428 24556 11480 24608
rect 11520 24556 11572 24608
rect 12532 24599 12584 24608
rect 12532 24565 12541 24599
rect 12541 24565 12575 24599
rect 12575 24565 12584 24599
rect 12532 24556 12584 24565
rect 13820 24556 13872 24608
rect 2663 24454 2715 24506
rect 2727 24454 2779 24506
rect 2791 24454 2843 24506
rect 2855 24454 2907 24506
rect 2919 24454 2971 24506
rect 6090 24454 6142 24506
rect 6154 24454 6206 24506
rect 6218 24454 6270 24506
rect 6282 24454 6334 24506
rect 6346 24454 6398 24506
rect 9517 24454 9569 24506
rect 9581 24454 9633 24506
rect 9645 24454 9697 24506
rect 9709 24454 9761 24506
rect 9773 24454 9825 24506
rect 12944 24454 12996 24506
rect 13008 24454 13060 24506
rect 13072 24454 13124 24506
rect 13136 24454 13188 24506
rect 13200 24454 13252 24506
rect 4896 24148 4948 24200
rect 7380 24352 7432 24404
rect 7472 24352 7524 24404
rect 6736 24284 6788 24336
rect 11244 24352 11296 24404
rect 11888 24352 11940 24404
rect 12164 24352 12216 24404
rect 8668 24216 8720 24268
rect 11428 24327 11480 24336
rect 11428 24293 11437 24327
rect 11437 24293 11471 24327
rect 11471 24293 11480 24327
rect 11428 24284 11480 24293
rect 11888 24216 11940 24268
rect 12532 24352 12584 24404
rect 13544 24352 13596 24404
rect 12624 24216 12676 24268
rect 13544 24216 13596 24268
rect 6368 24148 6420 24200
rect 6736 24148 6788 24200
rect 7104 24191 7156 24200
rect 7104 24157 7113 24191
rect 7113 24157 7147 24191
rect 7147 24157 7156 24191
rect 7104 24148 7156 24157
rect 7840 24191 7892 24200
rect 7840 24157 7849 24191
rect 7849 24157 7883 24191
rect 7883 24157 7892 24191
rect 7840 24148 7892 24157
rect 9128 24148 9180 24200
rect 9312 24148 9364 24200
rect 10784 24191 10836 24200
rect 10784 24157 10793 24191
rect 10793 24157 10827 24191
rect 10827 24157 10836 24191
rect 10784 24148 10836 24157
rect 756 24080 808 24132
rect 4988 24080 5040 24132
rect 8668 24080 8720 24132
rect 7564 24012 7616 24064
rect 13176 24123 13228 24132
rect 13176 24089 13185 24123
rect 13185 24089 13219 24123
rect 13219 24089 13228 24123
rect 13176 24080 13228 24089
rect 15108 24080 15160 24132
rect 11704 24012 11756 24064
rect 13268 24012 13320 24064
rect 13360 24012 13412 24064
rect 13728 24012 13780 24064
rect 4376 23910 4428 23962
rect 4440 23910 4492 23962
rect 4504 23910 4556 23962
rect 4568 23910 4620 23962
rect 4632 23910 4684 23962
rect 7803 23910 7855 23962
rect 7867 23910 7919 23962
rect 7931 23910 7983 23962
rect 7995 23910 8047 23962
rect 8059 23910 8111 23962
rect 11230 23910 11282 23962
rect 11294 23910 11346 23962
rect 11358 23910 11410 23962
rect 11422 23910 11474 23962
rect 11486 23910 11538 23962
rect 14657 23910 14709 23962
rect 14721 23910 14773 23962
rect 14785 23910 14837 23962
rect 14849 23910 14901 23962
rect 14913 23910 14965 23962
rect 3056 23672 3108 23724
rect 4896 23715 4948 23724
rect 4896 23681 4905 23715
rect 4905 23681 4939 23715
rect 4939 23681 4948 23715
rect 4896 23672 4948 23681
rect 5172 23715 5224 23724
rect 5172 23681 5179 23715
rect 5179 23681 5213 23715
rect 5213 23681 5224 23715
rect 5172 23672 5224 23681
rect 6828 23808 6880 23860
rect 8208 23851 8260 23860
rect 8208 23817 8217 23851
rect 8217 23817 8251 23851
rect 8251 23817 8260 23851
rect 8208 23808 8260 23817
rect 13176 23808 13228 23860
rect 10232 23740 10284 23792
rect 10784 23740 10836 23792
rect 12532 23740 12584 23792
rect 7288 23715 7340 23724
rect 7288 23681 7297 23715
rect 7297 23681 7331 23715
rect 7331 23681 7340 23715
rect 7288 23672 7340 23681
rect 7564 23715 7616 23724
rect 7564 23681 7573 23715
rect 7573 23681 7607 23715
rect 7607 23681 7616 23715
rect 7564 23672 7616 23681
rect 8852 23672 8904 23724
rect 12164 23715 12216 23724
rect 12164 23681 12173 23715
rect 12173 23681 12207 23715
rect 12207 23681 12216 23715
rect 12164 23672 12216 23681
rect 6000 23604 6052 23656
rect 6368 23647 6420 23656
rect 6368 23613 6377 23647
rect 6377 23613 6411 23647
rect 6411 23613 6420 23647
rect 6368 23604 6420 23613
rect 7380 23647 7432 23656
rect 7380 23613 7414 23647
rect 7414 23613 7432 23647
rect 7380 23604 7432 23613
rect 12072 23604 12124 23656
rect 12256 23604 12308 23656
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 12808 23647 12860 23656
rect 12808 23613 12817 23647
rect 12817 23613 12851 23647
rect 12851 23613 12860 23647
rect 12808 23604 12860 23613
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 13636 23647 13688 23656
rect 13636 23613 13670 23647
rect 13670 23613 13688 23647
rect 13636 23604 13688 23613
rect 13268 23579 13320 23588
rect 13268 23545 13277 23579
rect 13277 23545 13311 23579
rect 13311 23545 13320 23579
rect 13268 23536 13320 23545
rect 9220 23468 9272 23520
rect 10140 23511 10192 23520
rect 10140 23477 10149 23511
rect 10149 23477 10183 23511
rect 10183 23477 10192 23511
rect 10140 23468 10192 23477
rect 14188 23468 14240 23520
rect 2663 23366 2715 23418
rect 2727 23366 2779 23418
rect 2791 23366 2843 23418
rect 2855 23366 2907 23418
rect 2919 23366 2971 23418
rect 6090 23366 6142 23418
rect 6154 23366 6206 23418
rect 6218 23366 6270 23418
rect 6282 23366 6334 23418
rect 6346 23366 6398 23418
rect 9517 23366 9569 23418
rect 9581 23366 9633 23418
rect 9645 23366 9697 23418
rect 9709 23366 9761 23418
rect 9773 23366 9825 23418
rect 12944 23366 12996 23418
rect 13008 23366 13060 23418
rect 13072 23366 13124 23418
rect 13136 23366 13188 23418
rect 13200 23366 13252 23418
rect 5448 23264 5500 23316
rect 7196 23264 7248 23316
rect 7288 23264 7340 23316
rect 7472 23264 7524 23316
rect 12716 23264 12768 23316
rect 13268 23264 13320 23316
rect 9404 23128 9456 23180
rect 11704 23128 11756 23180
rect 11980 23128 12032 23180
rect 8852 23060 8904 23112
rect 10876 23060 10928 23112
rect 11152 23060 11204 23112
rect 12624 23103 12676 23112
rect 12624 23069 12631 23103
rect 12631 23069 12665 23103
rect 12665 23069 12676 23103
rect 12624 23060 12676 23069
rect 14372 23060 14424 23112
rect 756 22992 808 23044
rect 12992 22992 13044 23044
rect 10508 22924 10560 22976
rect 12624 22924 12676 22976
rect 12808 22924 12860 22976
rect 15108 22924 15160 22976
rect 4376 22822 4428 22874
rect 4440 22822 4492 22874
rect 4504 22822 4556 22874
rect 4568 22822 4620 22874
rect 4632 22822 4684 22874
rect 7803 22822 7855 22874
rect 7867 22822 7919 22874
rect 7931 22822 7983 22874
rect 7995 22822 8047 22874
rect 8059 22822 8111 22874
rect 11230 22822 11282 22874
rect 11294 22822 11346 22874
rect 11358 22822 11410 22874
rect 11422 22822 11474 22874
rect 11486 22822 11538 22874
rect 14657 22822 14709 22874
rect 14721 22822 14773 22874
rect 14785 22822 14837 22874
rect 14849 22822 14901 22874
rect 14913 22822 14965 22874
rect 1676 22720 1728 22772
rect 2320 22720 2372 22772
rect 10324 22720 10376 22772
rect 12992 22720 13044 22772
rect 756 22584 808 22636
rect 8392 22627 8444 22636
rect 8392 22593 8399 22627
rect 8399 22593 8433 22627
rect 8433 22593 8444 22627
rect 8392 22584 8444 22593
rect 9404 22584 9456 22636
rect 7748 22516 7800 22568
rect 10784 22516 10836 22568
rect 10876 22516 10928 22568
rect 12624 22584 12676 22636
rect 12716 22627 12768 22636
rect 12716 22593 12725 22627
rect 12725 22593 12759 22627
rect 12759 22593 12768 22627
rect 12716 22584 12768 22593
rect 9128 22423 9180 22432
rect 9128 22389 9137 22423
rect 9137 22389 9171 22423
rect 9171 22389 9180 22423
rect 9128 22380 9180 22389
rect 9404 22380 9456 22432
rect 13544 22720 13596 22772
rect 14280 22720 14332 22772
rect 14924 22720 14976 22772
rect 15292 22856 15344 22908
rect 15108 22788 15160 22840
rect 15476 22788 15528 22840
rect 15200 22720 15252 22772
rect 15384 22652 15436 22704
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 15936 22584 15988 22636
rect 13728 22516 13780 22568
rect 15660 22516 15712 22568
rect 14924 22448 14976 22500
rect 15292 22448 15344 22500
rect 13820 22423 13872 22432
rect 13820 22389 13829 22423
rect 13829 22389 13863 22423
rect 13863 22389 13872 22423
rect 13820 22380 13872 22389
rect 14372 22380 14424 22432
rect 15568 22380 15620 22432
rect 2663 22278 2715 22330
rect 2727 22278 2779 22330
rect 2791 22278 2843 22330
rect 2855 22278 2907 22330
rect 2919 22278 2971 22330
rect 6090 22278 6142 22330
rect 6154 22278 6206 22330
rect 6218 22278 6270 22330
rect 6282 22278 6334 22330
rect 6346 22278 6398 22330
rect 9517 22278 9569 22330
rect 9581 22278 9633 22330
rect 9645 22278 9697 22330
rect 9709 22278 9761 22330
rect 9773 22278 9825 22330
rect 12944 22278 12996 22330
rect 13008 22278 13060 22330
rect 13072 22278 13124 22330
rect 13136 22278 13188 22330
rect 13200 22278 13252 22330
rect 5172 22176 5224 22228
rect 5540 21972 5592 22024
rect 5908 21972 5960 22024
rect 6276 22015 6328 22024
rect 6276 21981 6285 22015
rect 6285 21981 6328 22015
rect 6276 21972 6328 21981
rect 7748 22176 7800 22228
rect 9036 22108 9088 22160
rect 7564 21972 7616 22024
rect 10784 22176 10836 22228
rect 11888 22176 11940 22228
rect 12900 22176 12952 22228
rect 13452 22176 13504 22228
rect 13636 22176 13688 22228
rect 14280 22219 14332 22228
rect 14280 22185 14289 22219
rect 14289 22185 14323 22219
rect 14323 22185 14332 22219
rect 14280 22176 14332 22185
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 10324 22108 10376 22160
rect 10140 22040 10192 22092
rect 10508 22040 10560 22092
rect 10968 22083 11020 22092
rect 10968 22049 10977 22083
rect 10977 22049 11011 22083
rect 11011 22049 11020 22083
rect 10968 22040 11020 22049
rect 7564 21836 7616 21888
rect 8392 21879 8444 21888
rect 8392 21845 8401 21879
rect 8401 21845 8435 21879
rect 8435 21845 8444 21879
rect 8392 21836 8444 21845
rect 10876 21972 10928 22024
rect 11980 21972 12032 22024
rect 12900 21972 12952 22024
rect 10324 21836 10376 21888
rect 10692 21836 10744 21888
rect 11612 21879 11664 21888
rect 11612 21845 11621 21879
rect 11621 21845 11655 21879
rect 11655 21845 11664 21879
rect 11612 21836 11664 21845
rect 12440 21836 12492 21888
rect 13452 21904 13504 21956
rect 14280 21972 14332 22024
rect 15844 21904 15896 21956
rect 13268 21836 13320 21888
rect 4376 21734 4428 21786
rect 4440 21734 4492 21786
rect 4504 21734 4556 21786
rect 4568 21734 4620 21786
rect 4632 21734 4684 21786
rect 7803 21734 7855 21786
rect 7867 21734 7919 21786
rect 7931 21734 7983 21786
rect 7995 21734 8047 21786
rect 8059 21734 8111 21786
rect 11230 21734 11282 21786
rect 11294 21734 11346 21786
rect 11358 21734 11410 21786
rect 11422 21734 11474 21786
rect 11486 21734 11538 21786
rect 14657 21734 14709 21786
rect 14721 21734 14773 21786
rect 14785 21734 14837 21786
rect 14849 21734 14901 21786
rect 14913 21734 14965 21786
rect 4988 21632 5040 21684
rect 756 21496 808 21548
rect 6828 21564 6880 21616
rect 7104 21564 7156 21616
rect 7472 21564 7524 21616
rect 7932 21564 7984 21616
rect 9864 21675 9916 21684
rect 9864 21641 9873 21675
rect 9873 21641 9907 21675
rect 9907 21641 9916 21675
rect 9864 21632 9916 21641
rect 12440 21632 12492 21684
rect 10692 21564 10744 21616
rect 13728 21632 13780 21684
rect 5908 21428 5960 21480
rect 7840 21428 7892 21480
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 8024 21428 8076 21437
rect 8392 21496 8444 21548
rect 9220 21539 9272 21548
rect 9220 21505 9229 21539
rect 9229 21505 9263 21539
rect 9263 21505 9272 21539
rect 9220 21496 9272 21505
rect 10876 21496 10928 21548
rect 12164 21539 12216 21548
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 8208 21292 8260 21344
rect 8760 21428 8812 21480
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 9128 21428 9180 21480
rect 12256 21428 12308 21480
rect 12900 21428 12952 21480
rect 13268 21471 13320 21480
rect 13268 21437 13277 21471
rect 13277 21437 13311 21471
rect 13311 21437 13320 21471
rect 13268 21428 13320 21437
rect 13636 21471 13688 21480
rect 13636 21437 13670 21471
rect 13670 21437 13688 21471
rect 13636 21428 13688 21437
rect 13820 21471 13872 21480
rect 13820 21437 13829 21471
rect 13829 21437 13863 21471
rect 13863 21437 13872 21471
rect 13820 21428 13872 21437
rect 14464 21428 14516 21480
rect 15936 21428 15988 21480
rect 10692 21292 10744 21344
rect 10968 21292 11020 21344
rect 12440 21292 12492 21344
rect 14280 21292 14332 21344
rect 2663 21190 2715 21242
rect 2727 21190 2779 21242
rect 2791 21190 2843 21242
rect 2855 21190 2907 21242
rect 2919 21190 2971 21242
rect 6090 21190 6142 21242
rect 6154 21190 6206 21242
rect 6218 21190 6270 21242
rect 6282 21190 6334 21242
rect 6346 21190 6398 21242
rect 9517 21190 9569 21242
rect 9581 21190 9633 21242
rect 9645 21190 9697 21242
rect 9709 21190 9761 21242
rect 9773 21190 9825 21242
rect 12944 21190 12996 21242
rect 13008 21190 13060 21242
rect 13072 21190 13124 21242
rect 13136 21190 13188 21242
rect 13200 21190 13252 21242
rect 3332 21131 3384 21140
rect 3332 21097 3341 21131
rect 3341 21097 3375 21131
rect 3375 21097 3384 21131
rect 3332 21088 3384 21097
rect 3240 21020 3292 21072
rect 6552 21020 6604 21072
rect 6736 21020 6788 21072
rect 6920 20952 6972 21004
rect 7380 21088 7432 21140
rect 7656 21088 7708 21140
rect 8024 21020 8076 21072
rect 7932 20952 7984 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 2504 20884 2556 20936
rect 6460 20884 6512 20936
rect 6552 20927 6604 20936
rect 6552 20893 6561 20927
rect 6561 20893 6595 20927
rect 6595 20893 6604 20927
rect 6552 20884 6604 20893
rect 7380 20927 7432 20936
rect 7380 20893 7414 20927
rect 7414 20893 7432 20927
rect 7380 20884 7432 20893
rect 7564 20927 7616 20936
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 8576 20884 8628 20936
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 8208 20816 8260 20868
rect 9680 20816 9732 20868
rect 6736 20748 6788 20800
rect 10508 20884 10560 20936
rect 10784 20791 10836 20800
rect 10784 20757 10793 20791
rect 10793 20757 10827 20791
rect 10827 20757 10836 20791
rect 10784 20748 10836 20757
rect 11152 20748 11204 20800
rect 13820 21088 13872 21140
rect 14096 21020 14148 21072
rect 11980 20952 12032 21004
rect 12256 20952 12308 21004
rect 12900 20927 12952 20936
rect 12164 20859 12216 20868
rect 12164 20825 12173 20859
rect 12173 20825 12207 20859
rect 12207 20825 12216 20859
rect 12164 20816 12216 20825
rect 12532 20859 12584 20868
rect 12532 20825 12541 20859
rect 12541 20825 12575 20859
rect 12575 20825 12584 20859
rect 12532 20816 12584 20825
rect 12900 20893 12925 20927
rect 12925 20893 12952 20927
rect 12900 20884 12952 20893
rect 13636 20748 13688 20800
rect 4376 20646 4428 20698
rect 4440 20646 4492 20698
rect 4504 20646 4556 20698
rect 4568 20646 4620 20698
rect 4632 20646 4684 20698
rect 7803 20646 7855 20698
rect 7867 20646 7919 20698
rect 7931 20646 7983 20698
rect 7995 20646 8047 20698
rect 8059 20646 8111 20698
rect 11230 20646 11282 20698
rect 11294 20646 11346 20698
rect 11358 20646 11410 20698
rect 11422 20646 11474 20698
rect 11486 20646 11538 20698
rect 14657 20646 14709 20698
rect 14721 20646 14773 20698
rect 14785 20646 14837 20698
rect 14849 20646 14901 20698
rect 14913 20646 14965 20698
rect 15936 20680 15988 20732
rect 4988 20544 5040 20596
rect 7932 20544 7984 20596
rect 4804 20383 4856 20392
rect 4804 20349 4813 20383
rect 4813 20349 4847 20383
rect 4847 20349 4856 20383
rect 4804 20340 4856 20349
rect 7288 20451 7340 20460
rect 7288 20417 7297 20451
rect 7297 20417 7331 20451
rect 7331 20417 7340 20451
rect 7288 20408 7340 20417
rect 9404 20476 9456 20528
rect 9680 20476 9732 20528
rect 10508 20476 10560 20528
rect 8392 20408 8444 20460
rect 7932 20340 7984 20392
rect 9404 20340 9456 20392
rect 11152 20544 11204 20596
rect 13912 20544 13964 20596
rect 15200 20544 15252 20596
rect 10784 20476 10836 20528
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 11612 20476 11664 20528
rect 7012 20204 7064 20256
rect 7196 20204 7248 20256
rect 7380 20247 7432 20256
rect 7380 20213 7389 20247
rect 7389 20213 7423 20247
rect 7423 20213 7432 20247
rect 7380 20204 7432 20213
rect 8576 20204 8628 20256
rect 9220 20247 9272 20256
rect 9220 20213 9229 20247
rect 9229 20213 9263 20247
rect 9263 20213 9272 20247
rect 9220 20204 9272 20213
rect 9312 20204 9364 20256
rect 11336 20272 11388 20324
rect 11612 20340 11664 20392
rect 12348 20408 12400 20460
rect 11060 20204 11112 20256
rect 11704 20204 11756 20256
rect 12256 20204 12308 20256
rect 12624 20204 12676 20256
rect 2663 20102 2715 20154
rect 2727 20102 2779 20154
rect 2791 20102 2843 20154
rect 2855 20102 2907 20154
rect 2919 20102 2971 20154
rect 6090 20102 6142 20154
rect 6154 20102 6206 20154
rect 6218 20102 6270 20154
rect 6282 20102 6334 20154
rect 6346 20102 6398 20154
rect 9517 20102 9569 20154
rect 9581 20102 9633 20154
rect 9645 20102 9697 20154
rect 9709 20102 9761 20154
rect 9773 20102 9825 20154
rect 12944 20102 12996 20154
rect 13008 20102 13060 20154
rect 13072 20102 13124 20154
rect 13136 20102 13188 20154
rect 13200 20102 13252 20154
rect 2412 20000 2464 20052
rect 5540 19932 5592 19984
rect 5816 19932 5868 19984
rect 756 19728 808 19780
rect 1124 19660 1176 19712
rect 7288 19932 7340 19984
rect 5816 19839 5868 19848
rect 5816 19805 5825 19839
rect 5825 19805 5859 19839
rect 5859 19805 5868 19839
rect 5816 19796 5868 19805
rect 6920 19796 6972 19848
rect 7104 19796 7156 19848
rect 7932 20000 7984 20052
rect 9220 20000 9272 20052
rect 8944 19907 8996 19916
rect 8944 19873 8953 19907
rect 8953 19873 8987 19907
rect 8987 19873 8996 19907
rect 8944 19864 8996 19873
rect 9862 19907 9914 19916
rect 9862 19873 9873 19907
rect 9873 19873 9907 19907
rect 9907 19873 9914 19907
rect 9862 19864 9914 19873
rect 10876 20000 10928 20052
rect 11796 20000 11848 20052
rect 12624 20000 12676 20052
rect 13820 20000 13872 20052
rect 8208 19796 8260 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 9956 19839 10008 19848
rect 12532 19932 12584 19984
rect 11336 19864 11388 19916
rect 12348 19864 12400 19916
rect 12808 19864 12860 19916
rect 13452 19864 13504 19916
rect 13636 19864 13688 19916
rect 9956 19805 9990 19839
rect 9990 19805 10008 19839
rect 9956 19796 10008 19805
rect 10692 19728 10744 19780
rect 13268 19839 13320 19848
rect 13268 19805 13277 19839
rect 13277 19805 13311 19839
rect 13311 19805 13320 19839
rect 13268 19796 13320 19805
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 9312 19660 9364 19712
rect 15200 19728 15252 19780
rect 15476 19728 15528 19780
rect 13820 19660 13872 19712
rect 4376 19558 4428 19610
rect 4440 19558 4492 19610
rect 4504 19558 4556 19610
rect 4568 19558 4620 19610
rect 4632 19558 4684 19610
rect 7803 19558 7855 19610
rect 7867 19558 7919 19610
rect 7931 19558 7983 19610
rect 7995 19558 8047 19610
rect 8059 19558 8111 19610
rect 11230 19558 11282 19610
rect 11294 19558 11346 19610
rect 11358 19558 11410 19610
rect 11422 19558 11474 19610
rect 11486 19558 11538 19610
rect 14657 19558 14709 19610
rect 14721 19558 14773 19610
rect 14785 19558 14837 19610
rect 14849 19558 14901 19610
rect 14913 19558 14965 19610
rect 7104 19456 7156 19508
rect 7196 19456 7248 19508
rect 6736 19388 6788 19440
rect 1492 19363 1544 19372
rect 1492 19329 1501 19363
rect 1501 19329 1535 19363
rect 1535 19329 1544 19363
rect 1492 19320 1544 19329
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 7748 19456 7800 19508
rect 9036 19456 9088 19508
rect 10876 19456 10928 19508
rect 11152 19456 11204 19508
rect 12532 19456 12584 19508
rect 7564 19320 7616 19372
rect 8208 19363 8260 19372
rect 8208 19329 8215 19363
rect 8215 19329 8249 19363
rect 8249 19329 8260 19363
rect 8208 19320 8260 19329
rect 10324 19320 10376 19372
rect 10600 19320 10652 19372
rect 7196 19263 7248 19315
rect 7380 19295 7432 19304
rect 7380 19261 7392 19295
rect 7392 19261 7426 19295
rect 7426 19261 7432 19295
rect 7380 19252 7432 19261
rect 10876 19320 10928 19372
rect 12256 19320 12308 19372
rect 3516 19184 3568 19236
rect 3608 19116 3660 19168
rect 5724 19116 5776 19168
rect 6000 19116 6052 19168
rect 7656 19116 7708 19168
rect 11704 19252 11756 19304
rect 13084 19320 13136 19372
rect 13268 19456 13320 19508
rect 14372 19499 14424 19508
rect 14372 19465 14381 19499
rect 14381 19465 14415 19499
rect 14415 19465 14424 19499
rect 14372 19456 14424 19465
rect 14464 19456 14516 19508
rect 14648 19456 14700 19508
rect 14464 19320 14516 19372
rect 9404 19184 9456 19236
rect 9956 19184 10008 19236
rect 10692 19184 10744 19236
rect 13820 19252 13872 19304
rect 8944 19159 8996 19168
rect 8944 19125 8953 19159
rect 8953 19125 8987 19159
rect 8987 19125 8996 19159
rect 8944 19116 8996 19125
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 12256 19116 12308 19168
rect 14096 19116 14148 19168
rect 2663 19014 2715 19066
rect 2727 19014 2779 19066
rect 2791 19014 2843 19066
rect 2855 19014 2907 19066
rect 2919 19014 2971 19066
rect 6090 19014 6142 19066
rect 6154 19014 6206 19066
rect 6218 19014 6270 19066
rect 6282 19014 6334 19066
rect 6346 19014 6398 19066
rect 9517 19014 9569 19066
rect 9581 19014 9633 19066
rect 9645 19014 9697 19066
rect 9709 19014 9761 19066
rect 9773 19014 9825 19066
rect 12944 19014 12996 19066
rect 13008 19014 13060 19066
rect 13072 19014 13124 19066
rect 13136 19014 13188 19066
rect 13200 19014 13252 19066
rect 3884 18912 3936 18964
rect 4712 18912 4764 18964
rect 8760 18912 8812 18964
rect 6920 18844 6972 18896
rect 7196 18844 7248 18896
rect 3976 18640 4028 18692
rect 5632 18708 5684 18760
rect 7656 18844 7708 18896
rect 7840 18844 7892 18896
rect 9680 18844 9732 18896
rect 5816 18640 5868 18692
rect 6000 18640 6052 18692
rect 7380 18708 7432 18760
rect 8576 18708 8628 18760
rect 9864 18751 9916 18760
rect 9864 18717 9873 18751
rect 9873 18717 9907 18751
rect 9907 18717 9916 18751
rect 9864 18708 9916 18717
rect 11980 18912 12032 18964
rect 14280 18912 14332 18964
rect 11612 18776 11664 18828
rect 11704 18776 11756 18828
rect 12256 18776 12308 18828
rect 10324 18640 10376 18692
rect 12348 18708 12400 18760
rect 12992 18708 13044 18760
rect 13820 18708 13872 18760
rect 14004 18708 14056 18760
rect 11612 18683 11664 18692
rect 11612 18649 11621 18683
rect 11621 18649 11655 18683
rect 11655 18649 11664 18683
rect 11612 18640 11664 18649
rect 12256 18640 12308 18692
rect 14556 18708 14608 18760
rect 6736 18572 6788 18624
rect 7104 18615 7156 18624
rect 7104 18581 7113 18615
rect 7113 18581 7147 18615
rect 7147 18581 7156 18615
rect 7104 18572 7156 18581
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 11152 18572 11204 18624
rect 11888 18572 11940 18624
rect 13544 18572 13596 18624
rect 13820 18572 13872 18624
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 4376 18470 4428 18522
rect 4440 18470 4492 18522
rect 4504 18470 4556 18522
rect 4568 18470 4620 18522
rect 4632 18470 4684 18522
rect 7803 18470 7855 18522
rect 7867 18470 7919 18522
rect 7931 18470 7983 18522
rect 7995 18470 8047 18522
rect 8059 18470 8111 18522
rect 11230 18470 11282 18522
rect 11294 18470 11346 18522
rect 11358 18470 11410 18522
rect 11422 18470 11474 18522
rect 11486 18470 11538 18522
rect 14657 18470 14709 18522
rect 14721 18470 14773 18522
rect 14785 18470 14837 18522
rect 14849 18470 14901 18522
rect 14913 18470 14965 18522
rect 6828 18411 6880 18420
rect 6828 18377 6837 18411
rect 6837 18377 6871 18411
rect 6871 18377 6880 18411
rect 6828 18368 6880 18377
rect 10876 18368 10928 18420
rect 11152 18368 11204 18420
rect 11888 18368 11940 18420
rect 756 18232 808 18284
rect 8668 18300 8720 18352
rect 3976 18232 4028 18284
rect 4252 18164 4304 18216
rect 4804 18207 4856 18216
rect 4804 18173 4813 18207
rect 4813 18173 4847 18207
rect 4847 18173 4856 18207
rect 4804 18164 4856 18173
rect 5816 18164 5868 18216
rect 6644 18164 6696 18216
rect 7472 18232 7524 18284
rect 7472 18096 7524 18148
rect 9588 18232 9640 18284
rect 9404 18164 9456 18216
rect 10140 18164 10192 18216
rect 11152 18275 11204 18284
rect 11152 18241 11161 18275
rect 11161 18241 11195 18275
rect 11195 18241 11204 18275
rect 11152 18232 11204 18241
rect 14096 18368 14148 18420
rect 14464 18411 14516 18420
rect 14464 18377 14473 18411
rect 14473 18377 14507 18411
rect 14507 18377 14516 18411
rect 14464 18368 14516 18377
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 12532 18164 12584 18216
rect 12716 18164 12768 18216
rect 12808 18207 12860 18216
rect 12808 18173 12817 18207
rect 12817 18173 12851 18207
rect 12851 18173 12860 18207
rect 12808 18164 12860 18173
rect 13636 18207 13688 18216
rect 13636 18173 13670 18207
rect 13670 18173 13688 18207
rect 13636 18164 13688 18173
rect 13268 18139 13320 18148
rect 13268 18105 13277 18139
rect 13277 18105 13311 18139
rect 13311 18105 13320 18139
rect 13268 18096 13320 18105
rect 6000 18028 6052 18080
rect 8576 18028 8628 18080
rect 9404 18028 9456 18080
rect 13360 18028 13412 18080
rect 13820 18028 13872 18080
rect 14464 18028 14516 18080
rect 2663 17926 2715 17978
rect 2727 17926 2779 17978
rect 2791 17926 2843 17978
rect 2855 17926 2907 17978
rect 2919 17926 2971 17978
rect 6090 17926 6142 17978
rect 6154 17926 6206 17978
rect 6218 17926 6270 17978
rect 6282 17926 6334 17978
rect 6346 17926 6398 17978
rect 9517 17926 9569 17978
rect 9581 17926 9633 17978
rect 9645 17926 9697 17978
rect 9709 17926 9761 17978
rect 9773 17926 9825 17978
rect 12944 17926 12996 17978
rect 13008 17926 13060 17978
rect 13072 17926 13124 17978
rect 13136 17926 13188 17978
rect 13200 17926 13252 17978
rect 7012 17824 7064 17876
rect 7564 17824 7616 17876
rect 8392 17824 8444 17876
rect 9220 17824 9272 17876
rect 5816 17756 5868 17808
rect 10692 17824 10744 17876
rect 11704 17824 11756 17876
rect 13268 17867 13320 17876
rect 13268 17833 13277 17867
rect 13277 17833 13311 17867
rect 13311 17833 13320 17867
rect 13268 17824 13320 17833
rect 13820 17867 13872 17876
rect 13820 17833 13829 17867
rect 13829 17833 13863 17867
rect 13863 17833 13872 17867
rect 13820 17824 13872 17833
rect 10876 17756 10928 17808
rect 8576 17688 8628 17740
rect 6000 17620 6052 17672
rect 756 17552 808 17604
rect 7104 17620 7156 17672
rect 9680 17663 9732 17672
rect 9680 17629 9687 17663
rect 9687 17629 9721 17663
rect 9721 17629 9732 17663
rect 9680 17620 9732 17629
rect 11704 17688 11756 17740
rect 12072 17688 12124 17740
rect 13544 17688 13596 17740
rect 14648 17688 14700 17740
rect 11428 17663 11480 17672
rect 11428 17629 11437 17663
rect 11437 17629 11471 17663
rect 11471 17629 11480 17663
rect 11428 17620 11480 17629
rect 11520 17620 11572 17672
rect 6460 17599 6485 17604
rect 6485 17599 6512 17604
rect 6460 17552 6512 17599
rect 12348 17552 12400 17604
rect 3608 17484 3660 17536
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 10692 17484 10744 17536
rect 10876 17484 10928 17536
rect 15200 17620 15252 17672
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 15200 17348 15252 17400
rect 15936 17348 15988 17400
rect 1676 17280 1728 17332
rect 7196 17280 7248 17332
rect 9312 17280 9364 17332
rect 1492 17187 1544 17196
rect 1492 17153 1501 17187
rect 1501 17153 1535 17187
rect 1535 17153 1544 17187
rect 1492 17144 1544 17153
rect 7012 17144 7064 17196
rect 11428 17212 11480 17264
rect 12624 17280 12676 17332
rect 13636 17280 13688 17332
rect 13912 17280 13964 17332
rect 15476 17280 15528 17332
rect 1400 17076 1452 17128
rect 1676 17076 1728 17128
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 7288 17076 7340 17085
rect 8208 17144 8260 17196
rect 9864 17144 9916 17196
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 13360 17144 13412 17196
rect 8300 17119 8352 17128
rect 8300 17085 8309 17119
rect 8309 17085 8343 17119
rect 8343 17085 8352 17119
rect 8300 17076 8352 17085
rect 9404 17076 9456 17128
rect 10048 16940 10100 16992
rect 10876 17076 10928 17128
rect 11244 17076 11296 17128
rect 12900 17076 12952 17128
rect 13452 17076 13504 17128
rect 10876 16940 10928 16992
rect 11704 16940 11756 16992
rect 12808 17008 12860 17060
rect 12716 16940 12768 16992
rect 13360 16940 13412 16992
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 1400 16736 1452 16788
rect 2504 16736 2556 16788
rect 6736 16736 6788 16788
rect 7104 16736 7156 16788
rect 8300 16736 8352 16788
rect 11796 16779 11848 16788
rect 11796 16745 11805 16779
rect 11805 16745 11839 16779
rect 11839 16745 11848 16779
rect 11796 16736 11848 16745
rect 12532 16736 12584 16788
rect 14372 16736 14424 16788
rect 8944 16668 8996 16720
rect 13912 16668 13964 16720
rect 6000 16600 6052 16652
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 10324 16600 10376 16652
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 11704 16600 11756 16652
rect 11796 16600 11848 16652
rect 11980 16600 12032 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 1768 16532 1820 16584
rect 8668 16532 8720 16584
rect 8852 16532 8904 16584
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 3884 16464 3936 16516
rect 5724 16464 5776 16516
rect 9588 16464 9640 16516
rect 1952 16396 2004 16448
rect 6552 16396 6604 16448
rect 7104 16396 7156 16448
rect 8484 16396 8536 16448
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 12900 16575 12952 16584
rect 12900 16541 12934 16575
rect 12934 16541 12952 16575
rect 12900 16532 12952 16541
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 13728 16464 13780 16516
rect 12440 16396 12492 16448
rect 12808 16396 12860 16448
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 6644 16192 6696 16244
rect 7104 16192 7156 16244
rect 8208 16124 8260 16176
rect 2044 16056 2096 16108
rect 6644 16056 6696 16108
rect 7564 16056 7616 16108
rect 11980 16192 12032 16244
rect 12532 16235 12584 16244
rect 12532 16201 12541 16235
rect 12541 16201 12575 16235
rect 12575 16201 12584 16235
rect 12532 16192 12584 16201
rect 10416 16167 10468 16176
rect 10416 16133 10425 16167
rect 10425 16133 10459 16167
rect 10459 16133 10468 16167
rect 10416 16124 10468 16133
rect 8944 16056 8996 16108
rect 10784 16056 10836 16108
rect 11060 16056 11112 16108
rect 13544 16056 13596 16108
rect 15476 16056 15528 16108
rect 15752 16056 15804 16108
rect 15936 16056 15988 16108
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 6736 15988 6788 16040
rect 6920 15920 6972 15972
rect 2412 15895 2464 15904
rect 2412 15861 2421 15895
rect 2421 15861 2455 15895
rect 2455 15861 2464 15895
rect 2412 15852 2464 15861
rect 9588 16031 9640 16040
rect 9588 15997 9622 16031
rect 9622 15997 9640 16031
rect 9588 15988 9640 15997
rect 9772 16031 9824 16040
rect 9772 15997 9781 16031
rect 9781 15997 9815 16031
rect 9815 15997 9824 16031
rect 9772 15988 9824 15997
rect 10416 15988 10468 16040
rect 11152 15988 11204 16040
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 12348 15988 12400 16040
rect 12808 15988 12860 16040
rect 12440 15920 12492 15972
rect 9128 15852 9180 15904
rect 11152 15852 11204 15904
rect 11612 15852 11664 15904
rect 12808 15852 12860 15904
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 5356 15648 5408 15700
rect 2320 15580 2372 15632
rect 6368 15580 6420 15632
rect 6920 15580 6972 15632
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 11060 15648 11112 15700
rect 11152 15648 11204 15700
rect 8576 15512 8628 15564
rect 756 15444 808 15496
rect 1584 15444 1636 15496
rect 1952 15487 2004 15496
rect 1952 15453 1961 15487
rect 1961 15453 1995 15487
rect 1995 15453 2004 15487
rect 1952 15444 2004 15453
rect 5080 15444 5132 15496
rect 9220 15487 9272 15496
rect 9220 15453 9227 15487
rect 9227 15453 9261 15487
rect 9261 15453 9272 15487
rect 9220 15444 9272 15453
rect 9772 15444 9824 15496
rect 13912 15648 13964 15700
rect 14372 15691 14424 15700
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 1768 15351 1820 15360
rect 1768 15317 1777 15351
rect 1777 15317 1811 15351
rect 1811 15317 1820 15351
rect 1768 15308 1820 15317
rect 5356 15308 5408 15360
rect 8300 15376 8352 15428
rect 10416 15376 10468 15428
rect 6460 15351 6512 15360
rect 6460 15317 6469 15351
rect 6469 15317 6503 15351
rect 6503 15317 6512 15351
rect 6460 15308 6512 15317
rect 8760 15308 8812 15360
rect 9220 15308 9272 15360
rect 14096 15512 14148 15564
rect 10784 15376 10836 15428
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 13084 15487 13136 15496
rect 13084 15453 13118 15487
rect 13118 15453 13136 15487
rect 13084 15444 13136 15453
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 14556 15444 14608 15496
rect 15752 15444 15804 15496
rect 10692 15308 10744 15360
rect 11612 15308 11664 15360
rect 11980 15308 12032 15360
rect 13084 15308 13136 15360
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 2412 15104 2464 15156
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 6736 15104 6788 15156
rect 8208 15104 8260 15156
rect 8300 15104 8352 15156
rect 1768 15036 1820 15088
rect 6368 15036 6420 15088
rect 12624 15104 12676 15156
rect 13268 15104 13320 15156
rect 6920 15011 6972 15020
rect 6920 14977 6929 15011
rect 6929 14977 6963 15011
rect 6963 14977 6972 15011
rect 6920 14968 6972 14977
rect 7104 14968 7156 15020
rect 6460 14900 6512 14952
rect 8576 14900 8628 14952
rect 9772 14943 9824 14952
rect 9772 14909 9781 14943
rect 9781 14909 9815 14943
rect 9815 14909 9824 14943
rect 9772 14900 9824 14909
rect 8392 14832 8444 14884
rect 9036 14832 9088 14884
rect 848 14764 900 14816
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 10048 14764 10100 14816
rect 10232 14764 10284 14816
rect 10784 14900 10836 14952
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 12072 15036 12124 15088
rect 11980 14968 12032 15020
rect 14188 15036 14240 15088
rect 12532 14900 12584 14952
rect 12716 14900 12768 14952
rect 11980 14875 12032 14884
rect 11980 14841 11989 14875
rect 11989 14841 12023 14875
rect 12023 14841 12032 14875
rect 11980 14832 12032 14841
rect 12072 14832 12124 14884
rect 12440 14832 12492 14884
rect 14556 14764 14608 14816
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 3792 14492 3844 14544
rect 5632 14492 5684 14544
rect 5080 14424 5132 14476
rect 5540 14424 5592 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 1676 14399 1728 14408
rect 1676 14365 1683 14399
rect 1683 14365 1717 14399
rect 1717 14365 1728 14399
rect 1676 14356 1728 14365
rect 1216 14288 1268 14340
rect 6920 14560 6972 14612
rect 7196 14492 7248 14544
rect 9128 14560 9180 14612
rect 9404 14560 9456 14612
rect 10784 14560 10836 14612
rect 9588 14492 9640 14544
rect 11520 14560 11572 14612
rect 11796 14560 11848 14612
rect 12164 14560 12216 14612
rect 13452 14560 13504 14612
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 7104 14220 7156 14272
rect 8852 14356 8904 14408
rect 9772 14356 9824 14408
rect 10508 14424 10560 14476
rect 10692 14424 10744 14476
rect 11152 14424 11204 14476
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 11980 14424 12032 14476
rect 10784 14356 10836 14408
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 12624 14467 12676 14476
rect 12624 14433 12633 14467
rect 12633 14433 12667 14467
rect 12667 14433 12676 14467
rect 12624 14424 12676 14433
rect 12348 14356 12400 14408
rect 13728 14356 13780 14408
rect 8300 14288 8352 14340
rect 8484 14288 8536 14340
rect 9588 14288 9640 14340
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 8852 14220 8904 14272
rect 11336 14220 11388 14272
rect 13820 14220 13872 14272
rect 14372 14220 14424 14272
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 848 14016 900 14068
rect 1952 14016 2004 14068
rect 2412 14016 2464 14068
rect 7104 14016 7156 14068
rect 7840 14016 7892 14068
rect 5816 13880 5868 13932
rect 9312 14016 9364 14068
rect 12072 14016 12124 14068
rect 12256 14016 12308 14068
rect 13636 14016 13688 14068
rect 15200 14016 15252 14068
rect 8852 13948 8904 14000
rect 9036 13991 9088 14000
rect 9036 13957 9045 13991
rect 9045 13957 9079 13991
rect 9079 13957 9088 13991
rect 9036 13948 9088 13957
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 10048 13948 10100 14000
rect 11060 13948 11112 14000
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 9772 13923 9824 13932
rect 9772 13889 9781 13923
rect 9781 13889 9815 13923
rect 9815 13889 9824 13923
rect 9772 13880 9824 13889
rect 10232 13880 10284 13932
rect 11704 13948 11756 14000
rect 11980 13948 12032 14000
rect 11796 13923 11848 13932
rect 11796 13889 11803 13923
rect 11803 13889 11837 13923
rect 11837 13889 11848 13923
rect 11796 13880 11848 13889
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 572 13812 624 13864
rect 4252 13812 4304 13864
rect 5448 13744 5500 13796
rect 5816 13744 5868 13796
rect 7196 13812 7248 13864
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 8300 13812 8352 13864
rect 8484 13812 8536 13864
rect 12624 13812 12676 13864
rect 7564 13787 7616 13796
rect 7564 13753 7573 13787
rect 7573 13753 7607 13787
rect 7607 13753 7616 13787
rect 7564 13744 7616 13753
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 7380 13676 7432 13728
rect 9036 13676 9088 13728
rect 10692 13676 10744 13728
rect 14004 13744 14056 13796
rect 14280 13744 14332 13796
rect 12532 13719 12584 13728
rect 12532 13685 12541 13719
rect 12541 13685 12575 13719
rect 12575 13685 12584 13719
rect 12532 13676 12584 13685
rect 13268 13676 13320 13728
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 5540 13336 5592 13388
rect 7564 13472 7616 13524
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 8484 13472 8536 13481
rect 9404 13472 9456 13524
rect 12532 13472 12584 13524
rect 12900 13472 12952 13524
rect 14280 13472 14332 13524
rect 14372 13515 14424 13524
rect 14372 13481 14381 13515
rect 14381 13481 14415 13515
rect 14415 13481 14424 13515
rect 14372 13472 14424 13481
rect 1952 13268 2004 13320
rect 5816 13268 5868 13320
rect 848 13132 900 13184
rect 10048 13336 10100 13388
rect 10324 13336 10376 13388
rect 11888 13336 11940 13388
rect 12256 13336 12308 13388
rect 13452 13404 13504 13456
rect 8576 13268 8628 13320
rect 8852 13268 8904 13320
rect 8208 13200 8260 13252
rect 11152 13268 11204 13320
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 14648 13336 14700 13388
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 15660 13268 15712 13320
rect 9404 13200 9456 13252
rect 9864 13132 9916 13184
rect 11244 13132 11296 13184
rect 13728 13132 13780 13184
rect 15844 13132 15896 13184
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 1584 12928 1636 12980
rect 4712 12928 4764 12980
rect 8576 12928 8628 12980
rect 11704 12928 11756 12980
rect 7104 12860 7156 12912
rect 6828 12792 6880 12844
rect 9404 12792 9456 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 10048 12792 10100 12844
rect 10784 12792 10836 12844
rect 11060 12792 11112 12844
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 12256 12792 12308 12844
rect 15200 12928 15252 12980
rect 12164 12724 12216 12776
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 12532 12724 12584 12776
rect 13636 12767 13688 12776
rect 13636 12733 13670 12767
rect 13670 12733 13688 12767
rect 13636 12724 13688 12733
rect 13268 12699 13320 12708
rect 13268 12665 13277 12699
rect 13277 12665 13311 12699
rect 13311 12665 13320 12699
rect 13268 12656 13320 12665
rect 14464 12699 14516 12708
rect 14464 12665 14473 12699
rect 14473 12665 14507 12699
rect 14507 12665 14516 12699
rect 14464 12656 14516 12665
rect 12440 12588 12492 12640
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 848 12384 900 12436
rect 9864 12384 9916 12436
rect 10692 12384 10744 12436
rect 8760 12316 8812 12368
rect 10416 12316 10468 12368
rect 10968 12316 11020 12368
rect 4896 12248 4948 12300
rect 5908 12248 5960 12300
rect 10232 12248 10284 12300
rect 10692 12248 10744 12300
rect 11888 12384 11940 12436
rect 12716 12384 12768 12436
rect 13452 12384 13504 12436
rect 13912 12427 13964 12436
rect 13912 12393 13921 12427
rect 13921 12393 13955 12427
rect 13955 12393 13964 12427
rect 13912 12384 13964 12393
rect 15936 12384 15988 12436
rect 14280 12316 14332 12368
rect 2412 12180 2464 12232
rect 9772 12180 9824 12232
rect 10600 12180 10652 12232
rect 12348 12180 12400 12232
rect 13268 12180 13320 12232
rect 13452 12180 13504 12232
rect 14188 12180 14240 12232
rect 15476 12180 15528 12232
rect 6644 12112 6696 12164
rect 9128 12112 9180 12164
rect 7564 12087 7616 12096
rect 7564 12053 7573 12087
rect 7573 12053 7607 12087
rect 7607 12053 7616 12087
rect 7564 12044 7616 12053
rect 9220 12044 9272 12096
rect 10324 12044 10376 12096
rect 11796 12044 11848 12096
rect 13820 12044 13872 12096
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 5264 11840 5316 11892
rect 12624 11840 12676 11892
rect 13636 11840 13688 11892
rect 13912 11840 13964 11892
rect 15568 11840 15620 11892
rect 5172 11777 5224 11824
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 5172 11772 5197 11777
rect 5197 11772 5224 11777
rect 7380 11704 7432 11756
rect 8852 11772 8904 11824
rect 9220 11772 9272 11824
rect 10048 11772 10100 11824
rect 10232 11815 10284 11824
rect 10232 11781 10241 11815
rect 10241 11781 10275 11815
rect 10275 11781 10284 11815
rect 10232 11772 10284 11781
rect 9772 11704 9824 11756
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 6828 11636 6880 11688
rect 7288 11636 7340 11688
rect 7472 11636 7524 11688
rect 1032 11568 1084 11620
rect 848 11500 900 11552
rect 6920 11500 6972 11552
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 7288 11500 7340 11552
rect 7472 11500 7524 11552
rect 8392 11500 8444 11552
rect 10692 11704 10744 11756
rect 11152 11636 11204 11688
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 13636 11747 13688 11756
rect 13636 11713 13670 11747
rect 13670 11713 13688 11747
rect 13636 11704 13688 11713
rect 13820 11747 13872 11756
rect 13820 11713 13829 11747
rect 13829 11713 13863 11747
rect 13863 11713 13872 11747
rect 13820 11704 13872 11713
rect 13268 11611 13320 11620
rect 13268 11577 13277 11611
rect 13277 11577 13311 11611
rect 13311 11577 13320 11611
rect 13268 11568 13320 11577
rect 12256 11500 12308 11552
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 4896 11160 4948 11212
rect 7472 11296 7524 11348
rect 8760 11296 8812 11348
rect 8852 11296 8904 11348
rect 9864 11296 9916 11348
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 10876 11296 10928 11348
rect 6828 11160 6880 11212
rect 6552 11092 6604 11144
rect 7472 11160 7524 11212
rect 11152 11228 11204 11280
rect 11244 11228 11296 11280
rect 13268 11296 13320 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 14464 11339 14516 11348
rect 14464 11305 14473 11339
rect 14473 11305 14507 11339
rect 14507 11305 14516 11339
rect 14464 11296 14516 11305
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 10232 11160 10284 11212
rect 11888 11160 11940 11212
rect 9312 11135 9364 11144
rect 9312 11101 9319 11135
rect 9319 11101 9353 11135
rect 9353 11101 9364 11135
rect 9312 11092 9364 11101
rect 2412 11024 2464 11076
rect 3884 11024 3936 11076
rect 4988 11024 5040 11076
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 6460 10956 6512 11008
rect 6644 10999 6696 11008
rect 6644 10965 6653 10999
rect 6653 10965 6687 10999
rect 6687 10965 6696 10999
rect 6644 10956 6696 10965
rect 6736 10956 6788 11008
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 8944 11024 8996 11076
rect 11060 11092 11112 11144
rect 11980 11092 12032 11144
rect 14648 11160 14700 11212
rect 10600 10956 10652 11008
rect 11612 11024 11664 11076
rect 14188 11092 14240 11144
rect 15108 11092 15160 11144
rect 12164 11024 12216 11076
rect 12716 10956 12768 11008
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 15844 10888 15896 10940
rect 1492 10752 1544 10804
rect 7012 10752 7064 10804
rect 7564 10752 7616 10804
rect 7748 10752 7800 10804
rect 10784 10752 10836 10804
rect 6736 10684 6788 10736
rect 11796 10684 11848 10736
rect 11980 10752 12032 10804
rect 12164 10752 12216 10804
rect 13820 10795 13872 10804
rect 13820 10761 13829 10795
rect 13829 10761 13863 10795
rect 13863 10761 13872 10795
rect 13820 10752 13872 10761
rect 6644 10616 6696 10668
rect 6460 10548 6512 10600
rect 6828 10548 6880 10600
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 8484 10616 8536 10668
rect 9312 10616 9364 10668
rect 12348 10616 12400 10668
rect 6920 10480 6972 10532
rect 4160 10412 4212 10464
rect 4252 10412 4304 10464
rect 6828 10412 6880 10464
rect 10692 10480 10744 10532
rect 11244 10480 11296 10532
rect 12164 10548 12216 10600
rect 14188 10659 14240 10668
rect 14188 10625 14197 10659
rect 14197 10625 14231 10659
rect 14231 10625 14240 10659
rect 14188 10616 14240 10625
rect 12716 10548 12768 10600
rect 7472 10412 7524 10464
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 11704 10412 11756 10464
rect 12440 10412 12492 10464
rect 15476 10412 15528 10464
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 7380 10208 7432 10260
rect 8392 10208 8444 10260
rect 10324 10208 10376 10260
rect 11060 10208 11112 10260
rect 12256 10208 12308 10260
rect 12624 10208 12676 10260
rect 12716 10208 12768 10260
rect 12992 10208 13044 10260
rect 13636 10208 13688 10260
rect 14004 10208 14056 10260
rect 3976 10140 4028 10192
rect 1032 10004 1084 10056
rect 2780 9936 2832 9988
rect 6460 10004 6512 10056
rect 9680 10072 9732 10124
rect 10232 10072 10284 10124
rect 10600 10072 10652 10124
rect 11244 10072 11296 10124
rect 11612 10072 11664 10124
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 12808 10072 12860 10124
rect 13452 10072 13504 10124
rect 8760 10004 8812 10056
rect 6644 9936 6696 9988
rect 9312 9936 9364 9988
rect 9496 9936 9548 9988
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 14280 9979 14332 9988
rect 14280 9945 14289 9979
rect 14289 9945 14323 9979
rect 14323 9945 14332 9979
rect 14280 9936 14332 9945
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 4160 9868 4212 9920
rect 10968 9868 11020 9920
rect 11612 9868 11664 9920
rect 11980 9868 12032 9920
rect 12256 9868 12308 9920
rect 12716 9868 12768 9920
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 2780 9707 2832 9716
rect 2780 9673 2789 9707
rect 2789 9673 2823 9707
rect 2823 9673 2832 9707
rect 2780 9664 2832 9673
rect 10416 9664 10468 9716
rect 10784 9664 10836 9716
rect 10968 9664 11020 9716
rect 13452 9664 13504 9716
rect 6552 9596 6604 9648
rect 7380 9596 7432 9648
rect 7656 9596 7708 9648
rect 11612 9596 11664 9648
rect 1768 9528 1820 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 6460 9571 6512 9580
rect 6460 9537 6469 9571
rect 6469 9537 6503 9571
rect 6503 9537 6512 9571
rect 6460 9528 6512 9537
rect 6920 9528 6972 9580
rect 7104 9528 7156 9580
rect 9496 9571 9548 9580
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 10600 9528 10652 9580
rect 12532 9528 12584 9580
rect 12716 9571 12768 9580
rect 12716 9537 12725 9571
rect 12725 9537 12759 9571
rect 12759 9537 12768 9571
rect 12716 9528 12768 9537
rect 8300 9460 8352 9512
rect 7472 9392 7524 9444
rect 8944 9392 8996 9444
rect 9864 9392 9916 9444
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 7840 9324 7892 9376
rect 10048 9460 10100 9512
rect 10876 9460 10928 9512
rect 11244 9460 11296 9512
rect 11428 9460 11480 9512
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 13820 9460 13872 9512
rect 10048 9324 10100 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 13360 9324 13412 9333
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 1124 9120 1176 9172
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 6460 9120 6512 9172
rect 6552 9120 6604 9172
rect 6644 9120 6696 9172
rect 8024 9120 8076 9172
rect 4896 8984 4948 9036
rect 8576 9052 8628 9104
rect 8944 9052 8996 9104
rect 7472 8984 7524 9036
rect 7656 8984 7708 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 8024 8984 8076 9036
rect 8484 8984 8536 9036
rect 10140 9120 10192 9172
rect 10508 9120 10560 9172
rect 11060 9120 11112 9172
rect 11336 9120 11388 9172
rect 13360 9120 13412 9172
rect 13452 9120 13504 9172
rect 9864 9027 9916 9036
rect 9864 8993 9873 9027
rect 9873 8993 9907 9027
rect 9907 8993 9916 9027
rect 9864 8984 9916 8993
rect 10324 8984 10376 9036
rect 10968 8984 11020 9036
rect 11796 9095 11848 9104
rect 11796 9061 11805 9095
rect 11805 9061 11839 9095
rect 11839 9061 11848 9095
rect 11796 9052 11848 9061
rect 13544 9052 13596 9104
rect 13636 8984 13688 9036
rect 1860 8848 1912 8900
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 8760 8916 8812 8968
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 9588 8916 9640 8968
rect 10140 8959 10192 8968
rect 10140 8925 10167 8959
rect 10167 8925 10192 8959
rect 10140 8916 10192 8925
rect 11244 8916 11296 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 15108 8916 15160 8968
rect 13360 8891 13412 8900
rect 13360 8857 13369 8891
rect 13369 8857 13403 8891
rect 13403 8857 13412 8891
rect 13360 8848 13412 8857
rect 13728 8891 13780 8900
rect 13728 8857 13737 8891
rect 13737 8857 13771 8891
rect 13771 8857 13780 8891
rect 13728 8848 13780 8857
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2412 8780 2464 8789
rect 5448 8780 5500 8832
rect 7472 8780 7524 8832
rect 9864 8780 9916 8832
rect 10048 8780 10100 8832
rect 11704 8780 11756 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 2412 8576 2464 8628
rect 6644 8576 6696 8628
rect 6920 8619 6972 8628
rect 6920 8585 6929 8619
rect 6929 8585 6963 8619
rect 6963 8585 6972 8619
rect 6920 8576 6972 8585
rect 7472 8576 7524 8628
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 9588 8576 9640 8628
rect 11612 8576 11664 8628
rect 11796 8576 11848 8628
rect 9864 8440 9916 8492
rect 10508 8483 10560 8492
rect 10508 8449 10542 8483
rect 10542 8449 10560 8483
rect 10508 8440 10560 8449
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 7196 8372 7248 8424
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 1676 8347 1728 8356
rect 1676 8313 1685 8347
rect 1685 8313 1719 8347
rect 1719 8313 1728 8347
rect 1676 8304 1728 8313
rect 7656 8304 7708 8356
rect 7932 8236 7984 8288
rect 8484 8236 8536 8288
rect 9772 8372 9824 8424
rect 12440 8508 12492 8560
rect 11888 8440 11940 8492
rect 12992 8576 13044 8628
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 12808 8508 12860 8560
rect 9864 8304 9916 8356
rect 10232 8304 10284 8356
rect 11336 8347 11388 8356
rect 11336 8313 11345 8347
rect 11345 8313 11379 8347
rect 11379 8313 11388 8347
rect 11336 8304 11388 8313
rect 11428 8304 11480 8356
rect 10876 8236 10928 8288
rect 11060 8236 11112 8288
rect 12624 8236 12676 8288
rect 12900 8236 12952 8288
rect 13820 8236 13872 8288
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 7656 8032 7708 8084
rect 7932 8032 7984 8084
rect 8760 8032 8812 8084
rect 11888 8032 11940 8084
rect 12348 8032 12400 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 13912 7964 13964 8016
rect 4896 7896 4948 7948
rect 1492 7803 1544 7812
rect 1492 7769 1501 7803
rect 1501 7769 1535 7803
rect 1535 7769 1544 7803
rect 1492 7760 1544 7769
rect 11520 7896 11572 7948
rect 6920 7760 6972 7812
rect 10876 7828 10928 7880
rect 11428 7828 11480 7880
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 12256 7828 12308 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 8392 7760 8444 7812
rect 12624 7760 12676 7812
rect 15108 7760 15160 7812
rect 848 7692 900 7744
rect 9404 7692 9456 7744
rect 13636 7692 13688 7744
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 5632 7488 5684 7540
rect 6552 7488 6604 7540
rect 10692 7488 10744 7540
rect 10968 7488 11020 7540
rect 11152 7488 11204 7540
rect 13176 7488 13228 7540
rect 13636 7488 13688 7540
rect 14372 7531 14424 7540
rect 14372 7497 14381 7531
rect 14381 7497 14415 7531
rect 14415 7497 14424 7531
rect 14372 7488 14424 7497
rect 13544 7420 13596 7472
rect 7012 7352 7064 7404
rect 9036 7352 9088 7404
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10692 7352 10744 7361
rect 11796 7395 11848 7404
rect 11796 7361 11803 7395
rect 11803 7361 11837 7395
rect 11837 7361 11848 7395
rect 11796 7352 11848 7361
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 14004 7420 14056 7472
rect 13912 7352 13964 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 6920 7284 6972 7336
rect 7656 7284 7708 7336
rect 10048 7284 10100 7336
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 10876 7284 10928 7336
rect 11060 7284 11112 7336
rect 13268 7284 13320 7336
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 9956 7148 10008 7200
rect 10784 7148 10836 7200
rect 11612 7148 11664 7200
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 1492 6944 1544 6996
rect 3240 6944 3292 6996
rect 8392 6944 8444 6996
rect 10140 6944 10192 6996
rect 11888 6944 11940 6996
rect 9404 6851 9456 6860
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 10324 6808 10376 6860
rect 10600 6808 10652 6860
rect 12072 6808 12124 6860
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 2412 6740 2464 6792
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 13544 6808 13596 6860
rect 15200 6808 15252 6860
rect 848 6604 900 6656
rect 11152 6604 11204 6656
rect 12716 6672 12768 6724
rect 13360 6672 13412 6724
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 13636 6715 13688 6724
rect 13636 6681 13645 6715
rect 13645 6681 13679 6715
rect 13679 6681 13688 6715
rect 13636 6672 13688 6681
rect 13820 6604 13872 6656
rect 15108 6672 15160 6724
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 2320 6400 2372 6452
rect 10048 6400 10100 6452
rect 11152 6400 11204 6452
rect 12716 6400 12768 6452
rect 14188 6400 14240 6452
rect 1584 6264 1636 6316
rect 5816 6264 5868 6316
rect 9036 6264 9088 6316
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 13360 6332 13412 6384
rect 14372 6332 14424 6384
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 12532 6307 12584 6316
rect 12532 6273 12566 6307
rect 12566 6273 12584 6307
rect 12532 6264 12584 6273
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 7656 6196 7708 6248
rect 9680 6239 9732 6248
rect 9680 6205 9689 6239
rect 9689 6205 9723 6239
rect 9723 6205 9732 6239
rect 9680 6196 9732 6205
rect 9864 6196 9916 6248
rect 10416 6239 10468 6248
rect 9956 6128 10008 6180
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 10876 6196 10928 6248
rect 12164 6171 12216 6180
rect 12164 6137 12173 6171
rect 12173 6137 12207 6171
rect 12207 6137 12216 6171
rect 12164 6128 12216 6137
rect 14740 6264 14792 6316
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 848 5856 900 5908
rect 8484 5899 8536 5908
rect 8484 5865 8493 5899
rect 8493 5865 8527 5899
rect 8527 5865 8536 5899
rect 8484 5856 8536 5865
rect 9312 5856 9364 5908
rect 12716 5856 12768 5908
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 4252 5720 4304 5772
rect 7656 5652 7708 5704
rect 14188 5788 14240 5840
rect 8208 5720 8260 5772
rect 8300 5652 8352 5704
rect 9772 5720 9824 5772
rect 10784 5720 10836 5772
rect 11980 5720 12032 5772
rect 12624 5652 12676 5704
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 9312 5584 9364 5636
rect 4712 5516 4764 5568
rect 9956 5516 10008 5568
rect 10876 5584 10928 5636
rect 13360 5652 13412 5704
rect 14004 5652 14056 5704
rect 13728 5627 13780 5636
rect 13728 5593 13737 5627
rect 13737 5593 13771 5627
rect 13771 5593 13780 5627
rect 13728 5584 13780 5593
rect 15108 5584 15160 5636
rect 12808 5516 12860 5568
rect 13912 5516 13964 5568
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 9864 5312 9916 5364
rect 10600 5312 10652 5364
rect 13544 5312 13596 5364
rect 2136 5244 2188 5296
rect 3608 5244 3660 5296
rect 7380 5176 7432 5228
rect 7656 5176 7708 5228
rect 848 4972 900 5024
rect 8392 5219 8444 5228
rect 8392 5185 8399 5219
rect 8399 5185 8433 5219
rect 8433 5185 8444 5219
rect 8392 5176 8444 5185
rect 9404 5176 9456 5228
rect 11980 5176 12032 5228
rect 12532 5176 12584 5228
rect 12716 5176 12768 5228
rect 9772 4972 9824 5024
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 3884 4768 3936 4820
rect 9404 4768 9456 4820
rect 12164 4768 12216 4820
rect 13452 4768 13504 4820
rect 11796 4700 11848 4752
rect 9864 4632 9916 4684
rect 756 4564 808 4616
rect 8668 4496 8720 4548
rect 12532 4564 12584 4616
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12952 4607
rect 12900 4564 12952 4573
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 11796 4088 11848 4140
rect 12532 4020 12584 4072
rect 13820 3884 13872 3936
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 9220 3680 9272 3732
rect 13360 3612 13412 3664
rect 12348 3544 12400 3596
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 14188 3476 14240 3485
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 13636 3043 13688 3052
rect 13636 3009 13645 3043
rect 13645 3009 13679 3043
rect 13679 3009 13688 3043
rect 13636 3000 13688 3009
rect 14372 3000 14424 3052
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
rect 5816 2091 5868 2100
rect 5816 2057 5825 2091
rect 5825 2057 5859 2091
rect 5859 2057 5868 2091
rect 5816 2048 5868 2057
rect 6552 2091 6604 2100
rect 6552 2057 6561 2091
rect 6561 2057 6595 2091
rect 6595 2057 6604 2091
rect 6552 2048 6604 2057
rect 4068 1980 4120 2032
rect 7656 2048 7708 2100
rect 8852 2048 8904 2100
rect 9956 2048 10008 2100
rect 11796 2048 11848 2100
rect 12440 2091 12492 2100
rect 12440 2057 12449 2091
rect 12449 2057 12483 2091
rect 12483 2057 12492 2091
rect 12440 2048 12492 2057
rect 14188 2091 14240 2100
rect 14188 2057 14197 2091
rect 14197 2057 14231 2091
rect 14231 2057 14240 2091
rect 14188 2048 14240 2057
rect 8944 1980 8996 2032
rect 11060 2023 11112 2032
rect 11060 1989 11069 2023
rect 11069 1989 11103 2023
rect 11103 1989 11112 2023
rect 11060 1980 11112 1989
rect 13452 1980 13504 2032
rect 1308 1912 1360 1964
rect 3056 1955 3108 1964
rect 3056 1921 3065 1955
rect 3065 1921 3099 1955
rect 3099 1921 3108 1955
rect 3056 1912 3108 1921
rect 5724 1955 5776 1964
rect 5724 1921 5733 1955
rect 5733 1921 5767 1955
rect 5767 1921 5776 1955
rect 5724 1912 5776 1921
rect 6460 1955 6512 1964
rect 6460 1921 6469 1955
rect 6469 1921 6503 1955
rect 6503 1921 6512 1955
rect 6460 1912 6512 1921
rect 7196 1955 7248 1964
rect 7196 1921 7205 1955
rect 7205 1921 7239 1955
rect 7239 1921 7248 1955
rect 7196 1912 7248 1921
rect 7932 1955 7984 1964
rect 7932 1921 7941 1955
rect 7941 1921 7975 1955
rect 7975 1921 7984 1955
rect 7932 1912 7984 1921
rect 8576 1955 8628 1964
rect 8576 1921 8585 1955
rect 8585 1921 8619 1955
rect 8619 1921 8628 1955
rect 8576 1912 8628 1921
rect 9312 1955 9364 1964
rect 9312 1921 9321 1955
rect 9321 1921 9355 1955
rect 9355 1921 9364 1955
rect 9312 1912 9364 1921
rect 10140 1955 10192 1964
rect 10140 1921 10149 1955
rect 10149 1921 10183 1955
rect 10183 1921 10192 1955
rect 10140 1912 10192 1921
rect 10876 1955 10928 1964
rect 10876 1921 10885 1955
rect 10885 1921 10919 1955
rect 10919 1921 10928 1955
rect 10876 1912 10928 1921
rect 11612 1955 11664 1964
rect 11612 1921 11621 1955
rect 11621 1921 11655 1955
rect 11655 1921 11664 1955
rect 11612 1912 11664 1921
rect 12348 1955 12400 1964
rect 12348 1921 12357 1955
rect 12357 1921 12391 1955
rect 12391 1921 12400 1955
rect 12348 1912 12400 1921
rect 13268 1912 13320 1964
rect 13728 1955 13780 1964
rect 13728 1921 13737 1955
rect 13737 1921 13771 1955
rect 13771 1921 13780 1955
rect 13728 1912 13780 1921
rect 11152 1844 11204 1896
rect 15200 1844 15252 1896
rect 15384 1844 15436 1896
rect 7380 1776 7432 1828
rect 2663 1606 2715 1658
rect 2727 1606 2779 1658
rect 2791 1606 2843 1658
rect 2855 1606 2907 1658
rect 2919 1606 2971 1658
rect 6090 1606 6142 1658
rect 6154 1606 6206 1658
rect 6218 1606 6270 1658
rect 6282 1606 6334 1658
rect 6346 1606 6398 1658
rect 9517 1606 9569 1658
rect 9581 1606 9633 1658
rect 9645 1606 9697 1658
rect 9709 1606 9761 1658
rect 9773 1606 9825 1658
rect 12944 1606 12996 1658
rect 13008 1606 13060 1658
rect 13072 1606 13124 1658
rect 13136 1606 13188 1658
rect 13200 1606 13252 1658
rect 5724 1504 5776 1556
rect 6460 1504 6512 1556
rect 7196 1504 7248 1556
rect 7932 1504 7984 1556
rect 8576 1504 8628 1556
rect 9312 1504 9364 1556
rect 10140 1504 10192 1556
rect 10876 1504 10928 1556
rect 11612 1504 11664 1556
rect 12348 1504 12400 1556
rect 13268 1504 13320 1556
rect 13452 1547 13504 1556
rect 13452 1513 13461 1547
rect 13461 1513 13495 1547
rect 13495 1513 13504 1547
rect 13452 1504 13504 1513
rect 13728 1547 13780 1556
rect 13728 1513 13737 1547
rect 13737 1513 13771 1547
rect 13771 1513 13780 1547
rect 13728 1504 13780 1513
rect 12532 1368 12584 1420
rect 2136 1343 2188 1352
rect 2136 1309 2145 1343
rect 2145 1309 2179 1343
rect 2179 1309 2188 1343
rect 2136 1300 2188 1309
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 4620 1343 4672 1352
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 5356 1343 5408 1352
rect 5356 1309 5365 1343
rect 5365 1309 5399 1343
rect 5399 1309 5408 1343
rect 5356 1300 5408 1309
rect 5724 1300 5776 1352
rect 6460 1300 6512 1352
rect 7196 1300 7248 1352
rect 8208 1343 8260 1352
rect 8208 1309 8217 1343
rect 8217 1309 8251 1343
rect 8251 1309 8260 1343
rect 8208 1300 8260 1309
rect 8668 1300 8720 1352
rect 9680 1343 9732 1352
rect 9680 1309 9689 1343
rect 9689 1309 9723 1343
rect 9723 1309 9732 1343
rect 9680 1300 9732 1309
rect 10140 1300 10192 1352
rect 10876 1300 10928 1352
rect 11612 1300 11664 1352
rect 12348 1300 12400 1352
rect 1584 1232 1636 1284
rect 4252 1232 4304 1284
rect 5172 1275 5224 1284
rect 5172 1241 5181 1275
rect 5181 1241 5215 1275
rect 5215 1241 5224 1275
rect 5172 1232 5224 1241
rect 13360 1343 13412 1352
rect 13360 1309 13369 1343
rect 13369 1309 13403 1343
rect 13403 1309 13412 1343
rect 13360 1300 13412 1309
rect 13912 1343 13964 1352
rect 13912 1309 13921 1343
rect 13921 1309 13955 1343
rect 13955 1309 13964 1343
rect 13912 1300 13964 1309
rect 14556 1300 14608 1352
rect 15292 1300 15344 1352
rect 15292 1164 15344 1216
rect 4376 1062 4428 1114
rect 4440 1062 4492 1114
rect 4504 1062 4556 1114
rect 4568 1062 4620 1114
rect 4632 1062 4684 1114
rect 7803 1062 7855 1114
rect 7867 1062 7919 1114
rect 7931 1062 7983 1114
rect 7995 1062 8047 1114
rect 8059 1062 8111 1114
rect 11230 1062 11282 1114
rect 11294 1062 11346 1114
rect 11358 1062 11410 1114
rect 11422 1062 11474 1114
rect 11486 1062 11538 1114
rect 14657 1062 14709 1114
rect 14721 1062 14773 1114
rect 14785 1062 14837 1114
rect 14849 1062 14901 1114
rect 14913 1062 14965 1114
<< metal2 >>
rect 570 44962 626 45000
rect 1306 44962 1362 45000
rect 2042 44962 2098 45000
rect 2778 44962 2834 45000
rect 570 44934 888 44962
rect 570 44840 626 44934
rect 860 43382 888 44934
rect 1306 44934 1624 44962
rect 1306 44840 1362 44934
rect 1596 43450 1624 44934
rect 2042 44934 2360 44962
rect 2042 44840 2098 44934
rect 2332 43450 2360 44934
rect 2778 44934 2912 44962
rect 2778 44840 2834 44934
rect 2884 43450 2912 44934
rect 3514 44840 3570 45000
rect 4250 44840 4306 45000
rect 4986 44962 5042 45000
rect 5722 44962 5778 45000
rect 6458 44962 6514 45000
rect 7194 44962 7250 45000
rect 7930 44962 7986 45000
rect 4986 44934 5304 44962
rect 4986 44840 5042 44934
rect 3528 43450 3556 44840
rect 4264 43450 4292 44840
rect 4376 43548 4684 43557
rect 4376 43546 4382 43548
rect 4438 43546 4462 43548
rect 4518 43546 4542 43548
rect 4598 43546 4622 43548
rect 4678 43546 4684 43548
rect 4438 43494 4440 43546
rect 4620 43494 4622 43546
rect 4376 43492 4382 43494
rect 4438 43492 4462 43494
rect 4518 43492 4542 43494
rect 4598 43492 4622 43494
rect 4678 43492 4684 43494
rect 4376 43483 4684 43492
rect 5276 43450 5304 44934
rect 5722 44934 5948 44962
rect 5722 44840 5778 44934
rect 5920 43450 5948 44934
rect 6458 44934 6776 44962
rect 6458 44840 6514 44934
rect 6748 43450 6776 44934
rect 7194 44934 7512 44962
rect 7194 44840 7250 44934
rect 7484 43450 7512 44934
rect 7930 44934 8248 44962
rect 7930 44840 7986 44934
rect 7803 43548 8111 43557
rect 7803 43546 7809 43548
rect 7865 43546 7889 43548
rect 7945 43546 7969 43548
rect 8025 43546 8049 43548
rect 8105 43546 8111 43548
rect 7865 43494 7867 43546
rect 8047 43494 8049 43546
rect 7803 43492 7809 43494
rect 7865 43492 7889 43494
rect 7945 43492 7969 43494
rect 8025 43492 8049 43494
rect 8105 43492 8111 43494
rect 7803 43483 8111 43492
rect 8220 43450 8248 44934
rect 8666 44840 8722 45000
rect 9402 44840 9458 45000
rect 10138 44962 10194 45000
rect 10138 44934 10456 44962
rect 10138 44840 10194 44934
rect 8680 43450 8708 44840
rect 9416 43450 9444 44840
rect 10428 43450 10456 44934
rect 10874 44840 10930 45000
rect 11610 44962 11666 45000
rect 11610 44934 11928 44962
rect 11610 44840 11666 44934
rect 10888 43450 10916 44840
rect 11230 43548 11538 43557
rect 11230 43546 11236 43548
rect 11292 43546 11316 43548
rect 11372 43546 11396 43548
rect 11452 43546 11476 43548
rect 11532 43546 11538 43548
rect 11292 43494 11294 43546
rect 11474 43494 11476 43546
rect 11230 43492 11236 43494
rect 11292 43492 11316 43494
rect 11372 43492 11396 43494
rect 11452 43492 11476 43494
rect 11532 43492 11538 43494
rect 11230 43483 11538 43492
rect 11900 43450 11928 44934
rect 12346 44840 12402 45000
rect 13082 44840 13138 45000
rect 13818 44840 13874 45000
rect 14554 44840 14610 45000
rect 15290 44840 15346 45000
rect 12360 43450 12388 44840
rect 13096 43450 13124 44840
rect 1584 43444 1636 43450
rect 1584 43386 1636 43392
rect 2320 43444 2372 43450
rect 2320 43386 2372 43392
rect 2872 43444 2924 43450
rect 2872 43386 2924 43392
rect 3516 43444 3568 43450
rect 3516 43386 3568 43392
rect 4252 43444 4304 43450
rect 4252 43386 4304 43392
rect 5264 43444 5316 43450
rect 5264 43386 5316 43392
rect 5908 43444 5960 43450
rect 5908 43386 5960 43392
rect 6736 43444 6788 43450
rect 6736 43386 6788 43392
rect 7472 43444 7524 43450
rect 7472 43386 7524 43392
rect 8208 43444 8260 43450
rect 8208 43386 8260 43392
rect 8668 43444 8720 43450
rect 8668 43386 8720 43392
rect 9404 43444 9456 43450
rect 9404 43386 9456 43392
rect 10416 43444 10468 43450
rect 10416 43386 10468 43392
rect 10876 43444 10928 43450
rect 10876 43386 10928 43392
rect 11888 43444 11940 43450
rect 11888 43386 11940 43392
rect 12348 43444 12400 43450
rect 12348 43386 12400 43392
rect 13084 43444 13136 43450
rect 13084 43386 13136 43392
rect 848 43376 900 43382
rect 848 43318 900 43324
rect 1768 43308 1820 43314
rect 1768 43250 1820 43256
rect 2136 43308 2188 43314
rect 2136 43250 2188 43256
rect 3056 43308 3108 43314
rect 3056 43250 3108 43256
rect 3240 43308 3292 43314
rect 3240 43250 3292 43256
rect 3792 43308 3844 43314
rect 3792 43250 3844 43256
rect 4436 43308 4488 43314
rect 4436 43250 4488 43256
rect 5080 43308 5132 43314
rect 5080 43250 5132 43256
rect 5816 43308 5868 43314
rect 5816 43250 5868 43256
rect 6644 43308 6696 43314
rect 6644 43250 6696 43256
rect 7288 43308 7340 43314
rect 7288 43250 7340 43256
rect 8116 43308 8168 43314
rect 8116 43250 8168 43256
rect 8944 43308 8996 43314
rect 8944 43250 8996 43256
rect 9220 43308 9272 43314
rect 9220 43250 9272 43256
rect 10232 43308 10284 43314
rect 10232 43250 10284 43256
rect 11612 43308 11664 43314
rect 11612 43250 11664 43256
rect 12072 43308 12124 43314
rect 12072 43250 12124 43256
rect 12532 43308 12584 43314
rect 12532 43250 12584 43256
rect 12808 43308 12860 43314
rect 12808 43250 12860 43256
rect 13728 43308 13780 43314
rect 13728 43250 13780 43256
rect 1032 42084 1084 42090
rect 1032 42026 1084 42032
rect 756 41132 808 41138
rect 756 41074 808 41080
rect 768 40905 796 41074
rect 754 40896 810 40905
rect 754 40831 810 40840
rect 756 40520 808 40526
rect 756 40462 808 40468
rect 768 40089 796 40462
rect 754 40080 810 40089
rect 754 40015 810 40024
rect 756 39432 808 39438
rect 756 39374 808 39380
rect 768 39273 796 39374
rect 754 39264 810 39273
rect 754 39199 810 39208
rect 756 37868 808 37874
rect 756 37810 808 37816
rect 768 37641 796 37810
rect 754 37632 810 37641
rect 754 37567 810 37576
rect 756 37188 808 37194
rect 756 37130 808 37136
rect 768 36825 796 37130
rect 754 36816 810 36825
rect 754 36751 810 36760
rect 756 36100 808 36106
rect 756 36042 808 36048
rect 768 36009 796 36042
rect 754 36000 810 36009
rect 754 35935 810 35944
rect 756 35692 808 35698
rect 756 35634 808 35640
rect 768 35193 796 35634
rect 754 35184 810 35193
rect 754 35119 810 35128
rect 756 33992 808 33998
rect 756 33934 808 33940
rect 768 33561 796 33934
rect 754 33552 810 33561
rect 754 33487 810 33496
rect 756 32904 808 32910
rect 756 32846 808 32852
rect 768 32745 796 32846
rect 754 32736 810 32745
rect 754 32671 810 32680
rect 756 32428 808 32434
rect 756 32370 808 32376
rect 768 31929 796 32370
rect 754 31920 810 31929
rect 754 31855 810 31864
rect 756 31340 808 31346
rect 756 31282 808 31288
rect 768 31113 796 31282
rect 754 31104 810 31113
rect 754 31039 810 31048
rect 756 29640 808 29646
rect 756 29582 808 29588
rect 768 29481 796 29582
rect 754 29472 810 29481
rect 754 29407 810 29416
rect 756 28076 808 28082
rect 756 28018 808 28024
rect 768 27849 796 28018
rect 754 27840 810 27849
rect 754 27775 810 27784
rect 756 27396 808 27402
rect 756 27338 808 27344
rect 768 27033 796 27338
rect 754 27024 810 27033
rect 754 26959 810 26968
rect 756 25832 808 25838
rect 756 25774 808 25780
rect 768 25401 796 25774
rect 754 25392 810 25401
rect 754 25327 810 25336
rect 756 24812 808 24818
rect 756 24754 808 24760
rect 768 24585 796 24754
rect 754 24576 810 24585
rect 754 24511 810 24520
rect 756 24132 808 24138
rect 756 24074 808 24080
rect 768 23769 796 24074
rect 754 23760 810 23769
rect 754 23695 810 23704
rect 756 23044 808 23050
rect 756 22986 808 22992
rect 768 22953 796 22986
rect 754 22944 810 22953
rect 754 22879 810 22888
rect 756 22636 808 22642
rect 756 22578 808 22584
rect 768 22137 796 22578
rect 754 22128 810 22137
rect 754 22063 810 22072
rect 756 21548 808 21554
rect 756 21490 808 21496
rect 768 21321 796 21490
rect 754 21312 810 21321
rect 754 21247 810 21256
rect 756 19780 808 19786
rect 756 19722 808 19728
rect 768 19689 796 19722
rect 754 19680 810 19689
rect 754 19615 810 19624
rect 756 18284 808 18290
rect 756 18226 808 18232
rect 768 18057 796 18226
rect 754 18048 810 18057
rect 754 17983 810 17992
rect 756 17604 808 17610
rect 756 17546 808 17552
rect 768 17241 796 17546
rect 754 17232 810 17241
rect 754 17167 810 17176
rect 754 15600 810 15609
rect 754 15535 810 15544
rect 768 15502 796 15535
rect 756 15496 808 15502
rect 756 15438 808 15444
rect 848 14816 900 14822
rect 846 14784 848 14793
rect 900 14784 902 14793
rect 846 14719 902 14728
rect 848 14068 900 14074
rect 848 14010 900 14016
rect 860 13977 888 14010
rect 846 13968 902 13977
rect 846 13903 902 13912
rect 572 13864 624 13870
rect 572 13806 624 13812
rect 584 160 612 13806
rect 848 13184 900 13190
rect 846 13152 848 13161
rect 900 13152 902 13161
rect 846 13087 902 13096
rect 848 12436 900 12442
rect 848 12378 900 12384
rect 860 12345 888 12378
rect 846 12336 902 12345
rect 846 12271 902 12280
rect 1044 11626 1072 42026
rect 1584 39296 1636 39302
rect 1584 39238 1636 39244
rect 1596 39098 1624 39238
rect 1584 39092 1636 39098
rect 1584 39034 1636 39040
rect 1400 38956 1452 38962
rect 1400 38898 1452 38904
rect 1412 38593 1440 38898
rect 1398 38584 1454 38593
rect 1398 38519 1454 38528
rect 1780 35834 1808 43250
rect 2148 42362 2176 43250
rect 2663 43004 2971 43013
rect 2663 43002 2669 43004
rect 2725 43002 2749 43004
rect 2805 43002 2829 43004
rect 2885 43002 2909 43004
rect 2965 43002 2971 43004
rect 2725 42950 2727 43002
rect 2907 42950 2909 43002
rect 2663 42948 2669 42950
rect 2725 42948 2749 42950
rect 2805 42948 2829 42950
rect 2885 42948 2909 42950
rect 2965 42948 2971 42950
rect 2663 42939 2971 42948
rect 2136 42356 2188 42362
rect 2136 42298 2188 42304
rect 2228 42220 2280 42226
rect 2228 42162 2280 42168
rect 1768 35828 1820 35834
rect 1768 35770 1820 35776
rect 1952 35692 2004 35698
rect 1952 35634 2004 35640
rect 1964 35290 1992 35634
rect 1952 35284 2004 35290
rect 1952 35226 2004 35232
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1412 34513 1440 34546
rect 1398 34504 1454 34513
rect 1398 34439 1454 34448
rect 2240 32570 2268 42162
rect 2663 41916 2971 41925
rect 2663 41914 2669 41916
rect 2725 41914 2749 41916
rect 2805 41914 2829 41916
rect 2885 41914 2909 41916
rect 2965 41914 2971 41916
rect 2725 41862 2727 41914
rect 2907 41862 2909 41914
rect 2663 41860 2669 41862
rect 2725 41860 2749 41862
rect 2805 41860 2829 41862
rect 2885 41860 2909 41862
rect 2965 41860 2971 41862
rect 2663 41851 2971 41860
rect 2663 40828 2971 40837
rect 2663 40826 2669 40828
rect 2725 40826 2749 40828
rect 2805 40826 2829 40828
rect 2885 40826 2909 40828
rect 2965 40826 2971 40828
rect 2725 40774 2727 40826
rect 2907 40774 2909 40826
rect 2663 40772 2669 40774
rect 2725 40772 2749 40774
rect 2805 40772 2829 40774
rect 2885 40772 2909 40774
rect 2965 40772 2971 40774
rect 2663 40763 2971 40772
rect 2663 39740 2971 39749
rect 2663 39738 2669 39740
rect 2725 39738 2749 39740
rect 2805 39738 2829 39740
rect 2885 39738 2909 39740
rect 2965 39738 2971 39740
rect 2725 39686 2727 39738
rect 2907 39686 2909 39738
rect 2663 39684 2669 39686
rect 2725 39684 2749 39686
rect 2805 39684 2829 39686
rect 2885 39684 2909 39686
rect 2965 39684 2971 39686
rect 2663 39675 2971 39684
rect 2663 38652 2971 38661
rect 2663 38650 2669 38652
rect 2725 38650 2749 38652
rect 2805 38650 2829 38652
rect 2885 38650 2909 38652
rect 2965 38650 2971 38652
rect 2725 38598 2727 38650
rect 2907 38598 2909 38650
rect 2663 38596 2669 38598
rect 2725 38596 2749 38598
rect 2805 38596 2829 38598
rect 2885 38596 2909 38598
rect 2965 38596 2971 38598
rect 2663 38587 2971 38596
rect 2663 37564 2971 37573
rect 2663 37562 2669 37564
rect 2725 37562 2749 37564
rect 2805 37562 2829 37564
rect 2885 37562 2909 37564
rect 2965 37562 2971 37564
rect 2725 37510 2727 37562
rect 2907 37510 2909 37562
rect 2663 37508 2669 37510
rect 2725 37508 2749 37510
rect 2805 37508 2829 37510
rect 2885 37508 2909 37510
rect 2965 37508 2971 37510
rect 2663 37499 2971 37508
rect 2663 36476 2971 36485
rect 2663 36474 2669 36476
rect 2725 36474 2749 36476
rect 2805 36474 2829 36476
rect 2885 36474 2909 36476
rect 2965 36474 2971 36476
rect 2725 36422 2727 36474
rect 2907 36422 2909 36474
rect 2663 36420 2669 36422
rect 2725 36420 2749 36422
rect 2805 36420 2829 36422
rect 2885 36420 2909 36422
rect 2965 36420 2971 36422
rect 2663 36411 2971 36420
rect 2663 35388 2971 35397
rect 2663 35386 2669 35388
rect 2725 35386 2749 35388
rect 2805 35386 2829 35388
rect 2885 35386 2909 35388
rect 2965 35386 2971 35388
rect 2725 35334 2727 35386
rect 2907 35334 2909 35386
rect 2663 35332 2669 35334
rect 2725 35332 2749 35334
rect 2805 35332 2829 35334
rect 2885 35332 2909 35334
rect 2965 35332 2971 35334
rect 2663 35323 2971 35332
rect 2663 34300 2971 34309
rect 2663 34298 2669 34300
rect 2725 34298 2749 34300
rect 2805 34298 2829 34300
rect 2885 34298 2909 34300
rect 2965 34298 2971 34300
rect 2725 34246 2727 34298
rect 2907 34246 2909 34298
rect 2663 34244 2669 34246
rect 2725 34244 2749 34246
rect 2805 34244 2829 34246
rect 2885 34244 2909 34246
rect 2965 34244 2971 34246
rect 2663 34235 2971 34244
rect 2663 33212 2971 33221
rect 2663 33210 2669 33212
rect 2725 33210 2749 33212
rect 2805 33210 2829 33212
rect 2885 33210 2909 33212
rect 2965 33210 2971 33212
rect 2725 33158 2727 33210
rect 2907 33158 2909 33210
rect 2663 33156 2669 33158
rect 2725 33156 2749 33158
rect 2805 33156 2829 33158
rect 2885 33156 2909 33158
rect 2965 33156 2971 33158
rect 2663 33147 2971 33156
rect 2228 32564 2280 32570
rect 2228 32506 2280 32512
rect 2228 32428 2280 32434
rect 2228 32370 2280 32376
rect 1860 32224 1912 32230
rect 1860 32166 1912 32172
rect 1872 31822 1900 32166
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 1216 31136 1268 31142
rect 1216 31078 1268 31084
rect 1228 28558 1256 31078
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 30297 1440 30670
rect 1398 30288 1454 30297
rect 1398 30223 1454 30232
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1412 28937 1440 29106
rect 1398 28928 1454 28937
rect 1398 28863 1454 28872
rect 1216 28552 1268 28558
rect 1216 28494 1268 28500
rect 1124 19712 1176 19718
rect 1124 19654 1176 19660
rect 1032 11620 1084 11626
rect 1032 11562 1084 11568
rect 848 11552 900 11558
rect 846 11520 848 11529
rect 900 11520 902 11529
rect 846 11455 902 11464
rect 1032 10056 1084 10062
rect 1032 9998 1084 10004
rect 1044 9897 1072 9998
rect 1030 9888 1086 9897
rect 1030 9823 1086 9832
rect 1136 9178 1164 19654
rect 1228 14346 1256 28494
rect 1400 28212 1452 28218
rect 1400 28154 1452 28160
rect 1412 21434 1440 28154
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1596 26314 1624 27270
rect 1492 26308 1544 26314
rect 1492 26250 1544 26256
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1504 26217 1532 26250
rect 1490 26208 1546 26217
rect 1490 26143 1546 26152
rect 1412 21406 1532 21434
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20641 1440 20878
rect 1398 20632 1454 20641
rect 1398 20567 1454 20576
rect 1504 20482 1532 21406
rect 1412 20454 1532 20482
rect 1412 17134 1440 20454
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1504 19281 1532 19314
rect 1490 19272 1546 19281
rect 1490 19207 1546 19216
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1412 16590 1440 16730
rect 1400 16584 1452 16590
rect 1504 16561 1532 17138
rect 1400 16526 1452 16532
rect 1490 16552 1546 16561
rect 1412 16046 1440 16526
rect 1490 16487 1546 16496
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 14414 1440 15982
rect 1596 15502 1624 26250
rect 1674 23216 1730 23225
rect 1674 23151 1730 23160
rect 1688 22778 1716 23151
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 1674 19272 1730 19281
rect 1674 19207 1730 19216
rect 1688 17338 1716 19207
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1676 17128 1728 17134
rect 1676 17070 1728 17076
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1216 14340 1268 14346
rect 1216 14282 1268 14288
rect 1412 12782 1440 14350
rect 1596 12986 1624 15438
rect 1688 14414 1716 17070
rect 1780 16590 1808 29446
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1780 15094 1808 15302
rect 1768 15088 1820 15094
rect 1768 15030 1820 15036
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 9518 1440 12718
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 10810 1532 11698
rect 1584 11008 1636 11014
rect 1582 10976 1584 10985
rect 1636 10976 1638 10985
rect 1582 10911 1638 10920
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9625 1624 9862
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 1766 9616 1822 9625
rect 1766 9551 1768 9560
rect 1820 9551 1822 9560
rect 1768 9522 1820 9528
rect 1400 9512 1452 9518
rect 1872 9489 1900 31758
rect 2240 31346 2268 32370
rect 2663 32124 2971 32133
rect 2663 32122 2669 32124
rect 2725 32122 2749 32124
rect 2805 32122 2829 32124
rect 2885 32122 2909 32124
rect 2965 32122 2971 32124
rect 2725 32070 2727 32122
rect 2907 32070 2909 32122
rect 2663 32068 2669 32070
rect 2725 32068 2749 32070
rect 2805 32068 2829 32070
rect 2885 32068 2909 32070
rect 2965 32068 2971 32070
rect 2663 32059 2971 32068
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 2663 31036 2971 31045
rect 2663 31034 2669 31036
rect 2725 31034 2749 31036
rect 2805 31034 2829 31036
rect 2885 31034 2909 31036
rect 2965 31034 2971 31036
rect 2725 30982 2727 31034
rect 2907 30982 2909 31034
rect 2663 30980 2669 30982
rect 2725 30980 2749 30982
rect 2805 30980 2829 30982
rect 2885 30980 2909 30982
rect 2965 30980 2971 30982
rect 2663 30971 2971 30980
rect 2663 29948 2971 29957
rect 2663 29946 2669 29948
rect 2725 29946 2749 29948
rect 2805 29946 2829 29948
rect 2885 29946 2909 29948
rect 2965 29946 2971 29948
rect 2725 29894 2727 29946
rect 2907 29894 2909 29946
rect 2663 29892 2669 29894
rect 2725 29892 2749 29894
rect 2805 29892 2829 29894
rect 2885 29892 2909 29894
rect 2965 29892 2971 29894
rect 2663 29883 2971 29892
rect 2412 29164 2464 29170
rect 2412 29106 2464 29112
rect 1952 29028 2004 29034
rect 1952 28970 2004 28976
rect 1964 20369 1992 28970
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 1950 20360 2006 20369
rect 1950 20295 2006 20304
rect 1964 16574 1992 20295
rect 1964 16546 2084 16574
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 15502 1992 16390
rect 2056 16114 2084 16546
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2332 15638 2360 22714
rect 2424 20058 2452 29106
rect 2663 28860 2971 28869
rect 2663 28858 2669 28860
rect 2725 28858 2749 28860
rect 2805 28858 2829 28860
rect 2885 28858 2909 28860
rect 2965 28858 2971 28860
rect 2725 28806 2727 28858
rect 2907 28806 2909 28858
rect 2663 28804 2669 28806
rect 2725 28804 2749 28806
rect 2805 28804 2829 28806
rect 2885 28804 2909 28806
rect 2965 28804 2971 28806
rect 2663 28795 2971 28804
rect 2663 27772 2971 27781
rect 2663 27770 2669 27772
rect 2725 27770 2749 27772
rect 2805 27770 2829 27772
rect 2885 27770 2909 27772
rect 2965 27770 2971 27772
rect 2725 27718 2727 27770
rect 2907 27718 2909 27770
rect 2663 27716 2669 27718
rect 2725 27716 2749 27718
rect 2805 27716 2829 27718
rect 2885 27716 2909 27718
rect 2965 27716 2971 27718
rect 2663 27707 2971 27716
rect 3068 27130 3096 43250
rect 3252 42906 3280 43250
rect 3804 42906 3832 43250
rect 4448 42906 4476 43250
rect 5092 42906 5120 43250
rect 5828 42906 5856 43250
rect 6090 43004 6398 43013
rect 6090 43002 6096 43004
rect 6152 43002 6176 43004
rect 6232 43002 6256 43004
rect 6312 43002 6336 43004
rect 6392 43002 6398 43004
rect 6152 42950 6154 43002
rect 6334 42950 6336 43002
rect 6090 42948 6096 42950
rect 6152 42948 6176 42950
rect 6232 42948 6256 42950
rect 6312 42948 6336 42950
rect 6392 42948 6398 42950
rect 6090 42939 6398 42948
rect 6656 42906 6684 43250
rect 7300 42906 7328 43250
rect 8128 42906 8156 43250
rect 8956 42906 8984 43250
rect 9232 42906 9260 43250
rect 9517 43004 9825 43013
rect 9517 43002 9523 43004
rect 9579 43002 9603 43004
rect 9659 43002 9683 43004
rect 9739 43002 9763 43004
rect 9819 43002 9825 43004
rect 9579 42950 9581 43002
rect 9761 42950 9763 43002
rect 9517 42948 9523 42950
rect 9579 42948 9603 42950
rect 9659 42948 9683 42950
rect 9739 42948 9763 42950
rect 9819 42948 9825 42950
rect 9517 42939 9825 42948
rect 10244 42906 10272 43250
rect 11624 42906 11652 43250
rect 12084 42906 12112 43250
rect 12544 42906 12572 43250
rect 12820 42906 12848 43250
rect 12944 43004 13252 43013
rect 12944 43002 12950 43004
rect 13006 43002 13030 43004
rect 13086 43002 13110 43004
rect 13166 43002 13190 43004
rect 13246 43002 13252 43004
rect 13006 42950 13008 43002
rect 13188 42950 13190 43002
rect 12944 42948 12950 42950
rect 13006 42948 13030 42950
rect 13086 42948 13110 42950
rect 13166 42948 13190 42950
rect 13246 42948 13252 42950
rect 12944 42939 13252 42948
rect 3240 42900 3292 42906
rect 3240 42842 3292 42848
rect 3792 42900 3844 42906
rect 3792 42842 3844 42848
rect 4436 42900 4488 42906
rect 4436 42842 4488 42848
rect 5080 42900 5132 42906
rect 5080 42842 5132 42848
rect 5816 42900 5868 42906
rect 5816 42842 5868 42848
rect 6644 42900 6696 42906
rect 6644 42842 6696 42848
rect 7288 42900 7340 42906
rect 7288 42842 7340 42848
rect 8116 42900 8168 42906
rect 8116 42842 8168 42848
rect 8944 42900 8996 42906
rect 8944 42842 8996 42848
rect 9220 42900 9272 42906
rect 9220 42842 9272 42848
rect 10232 42900 10284 42906
rect 10232 42842 10284 42848
rect 11612 42900 11664 42906
rect 11612 42842 11664 42848
rect 12072 42900 12124 42906
rect 12072 42842 12124 42848
rect 12532 42900 12584 42906
rect 12532 42842 12584 42848
rect 12808 42900 12860 42906
rect 12808 42842 12860 42848
rect 3792 42764 3844 42770
rect 3792 42706 3844 42712
rect 3516 42696 3568 42702
rect 3516 42638 3568 42644
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 3056 26988 3108 26994
rect 3056 26930 3108 26936
rect 2663 26684 2971 26693
rect 2663 26682 2669 26684
rect 2725 26682 2749 26684
rect 2805 26682 2829 26684
rect 2885 26682 2909 26684
rect 2965 26682 2971 26684
rect 2725 26630 2727 26682
rect 2907 26630 2909 26682
rect 2663 26628 2669 26630
rect 2725 26628 2749 26630
rect 2805 26628 2829 26630
rect 2885 26628 2909 26630
rect 2965 26628 2971 26630
rect 2663 26619 2971 26628
rect 3068 26586 3096 26930
rect 3056 26580 3108 26586
rect 3056 26522 3108 26528
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 2663 25596 2971 25605
rect 2663 25594 2669 25596
rect 2725 25594 2749 25596
rect 2805 25594 2829 25596
rect 2885 25594 2909 25596
rect 2965 25594 2971 25596
rect 2725 25542 2727 25594
rect 2907 25542 2909 25594
rect 2663 25540 2669 25542
rect 2725 25540 2749 25542
rect 2805 25540 2829 25542
rect 2885 25540 2909 25542
rect 2965 25540 2971 25542
rect 2663 25531 2971 25540
rect 2663 24508 2971 24517
rect 2663 24506 2669 24508
rect 2725 24506 2749 24508
rect 2805 24506 2829 24508
rect 2885 24506 2909 24508
rect 2965 24506 2971 24508
rect 2725 24454 2727 24506
rect 2907 24454 2909 24506
rect 2663 24452 2669 24454
rect 2725 24452 2749 24454
rect 2805 24452 2829 24454
rect 2885 24452 2909 24454
rect 2965 24452 2971 24454
rect 2663 24443 2971 24452
rect 3068 23730 3096 26318
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 2663 23420 2971 23429
rect 2663 23418 2669 23420
rect 2725 23418 2749 23420
rect 2805 23418 2829 23420
rect 2885 23418 2909 23420
rect 2965 23418 2971 23420
rect 2725 23366 2727 23418
rect 2907 23366 2909 23418
rect 2663 23364 2669 23366
rect 2725 23364 2749 23366
rect 2805 23364 2829 23366
rect 2885 23364 2909 23366
rect 2965 23364 2971 23366
rect 2663 23355 2971 23364
rect 2663 22332 2971 22341
rect 2663 22330 2669 22332
rect 2725 22330 2749 22332
rect 2805 22330 2829 22332
rect 2885 22330 2909 22332
rect 2965 22330 2971 22332
rect 2725 22278 2727 22330
rect 2907 22278 2909 22330
rect 2663 22276 2669 22278
rect 2725 22276 2749 22278
rect 2805 22276 2829 22278
rect 2885 22276 2909 22278
rect 2965 22276 2971 22278
rect 2663 22267 2971 22276
rect 3528 22094 3556 42638
rect 3608 33856 3660 33862
rect 3608 33798 3660 33804
rect 3344 22066 3556 22094
rect 2663 21244 2971 21253
rect 2663 21242 2669 21244
rect 2725 21242 2749 21244
rect 2805 21242 2829 21244
rect 2885 21242 2909 21244
rect 2965 21242 2971 21244
rect 2725 21190 2727 21242
rect 2907 21190 2909 21242
rect 2663 21188 2669 21190
rect 2725 21188 2749 21190
rect 2805 21188 2829 21190
rect 2885 21188 2909 21190
rect 2965 21188 2971 21190
rect 2663 21179 2971 21188
rect 3344 21146 3372 22066
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2424 16574 2452 19994
rect 2516 16794 2544 20878
rect 2663 20156 2971 20165
rect 2663 20154 2669 20156
rect 2725 20154 2749 20156
rect 2805 20154 2829 20156
rect 2885 20154 2909 20156
rect 2965 20154 2971 20156
rect 2725 20102 2727 20154
rect 2907 20102 2909 20154
rect 2663 20100 2669 20102
rect 2725 20100 2749 20102
rect 2805 20100 2829 20102
rect 2885 20100 2909 20102
rect 2965 20100 2971 20102
rect 2663 20091 2971 20100
rect 2663 19068 2971 19077
rect 2663 19066 2669 19068
rect 2725 19066 2749 19068
rect 2805 19066 2829 19068
rect 2885 19066 2909 19068
rect 2965 19066 2971 19068
rect 2725 19014 2727 19066
rect 2907 19014 2909 19066
rect 2663 19012 2669 19014
rect 2725 19012 2749 19014
rect 2805 19012 2829 19014
rect 2885 19012 2909 19014
rect 2965 19012 2971 19014
rect 2663 19003 2971 19012
rect 2663 17980 2971 17989
rect 2663 17978 2669 17980
rect 2725 17978 2749 17980
rect 2805 17978 2829 17980
rect 2885 17978 2909 17980
rect 2965 17978 2971 17980
rect 2725 17926 2727 17978
rect 2907 17926 2909 17978
rect 2663 17924 2669 17926
rect 2725 17924 2749 17926
rect 2805 17924 2829 17926
rect 2885 17924 2909 17926
rect 2965 17924 2971 17926
rect 2663 17915 2971 17924
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2424 16546 2544 16574
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2320 15632 2372 15638
rect 2320 15574 2372 15580
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 2424 15162 2452 15846
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14074 1992 14758
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2424 14074 2452 14214
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13326 1992 13670
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 12238 2452 12582
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2424 10266 2452 11018
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 1400 9454 1452 9460
rect 1858 9480 1914 9489
rect 1124 9172 1176 9178
rect 1124 9114 1176 9120
rect 1412 8974 1440 9454
rect 1858 9415 1914 9424
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 848 7744 900 7750
rect 848 7686 900 7692
rect 860 7449 888 7686
rect 846 7440 902 7449
rect 846 7375 902 7384
rect 1412 7342 1440 8910
rect 1872 8906 1900 9415
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2424 8634 2452 8774
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1688 8265 1716 8298
rect 1674 8256 1730 8265
rect 1674 8191 1730 8200
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 848 6656 900 6662
rect 846 6624 848 6633
rect 900 6624 902 6633
rect 846 6559 902 6568
rect 1412 6338 1440 7278
rect 1504 7002 1532 7754
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 2424 6798 2452 7142
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2332 6458 2360 6734
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 1412 6322 1624 6338
rect 1412 6316 1636 6322
rect 1412 6310 1584 6316
rect 1584 6258 1636 6264
rect 848 5908 900 5914
rect 848 5850 900 5856
rect 860 5817 888 5850
rect 846 5808 902 5817
rect 846 5743 902 5752
rect 848 5024 900 5030
rect 846 4992 848 5001
rect 900 4992 902 5001
rect 846 4927 902 4936
rect 756 4616 808 4622
rect 756 4558 808 4564
rect 768 4185 796 4558
rect 754 4176 810 4185
rect 754 4111 810 4120
rect 1308 1964 1360 1970
rect 1308 1906 1360 1912
rect 1320 160 1348 1906
rect 1596 1290 1624 6258
rect 2516 5681 2544 16546
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2792 9722 2820 9930
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 3252 7002 3280 21014
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3528 18873 3556 19178
rect 3620 19174 3648 33798
rect 3804 19334 3832 42706
rect 4068 42696 4120 42702
rect 4068 42638 4120 42644
rect 5080 42696 5132 42702
rect 5080 42638 5132 42644
rect 7288 42696 7340 42702
rect 7288 42638 7340 42644
rect 7472 42696 7524 42702
rect 7472 42638 7524 42644
rect 9404 42696 9456 42702
rect 9404 42638 9456 42644
rect 10968 42696 11020 42702
rect 10968 42638 11020 42644
rect 11704 42696 11756 42702
rect 12440 42696 12492 42702
rect 11704 42638 11756 42644
rect 12438 42664 12440 42673
rect 12492 42664 12494 42673
rect 3976 42560 4028 42566
rect 3976 42502 4028 42508
rect 3884 42288 3936 42294
rect 3884 42230 3936 42236
rect 3712 19306 3832 19334
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3514 18864 3570 18873
rect 3514 18799 3570 18808
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2148 5302 2176 5510
rect 3620 5302 3648 17478
rect 3712 14532 3740 19306
rect 3896 18970 3924 42230
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 3988 18816 4016 42502
rect 4080 42362 4108 42638
rect 4804 42628 4856 42634
rect 4804 42570 4856 42576
rect 4376 42460 4684 42469
rect 4376 42458 4382 42460
rect 4438 42458 4462 42460
rect 4518 42458 4542 42460
rect 4598 42458 4622 42460
rect 4678 42458 4684 42460
rect 4438 42406 4440 42458
rect 4620 42406 4622 42458
rect 4376 42404 4382 42406
rect 4438 42404 4462 42406
rect 4518 42404 4542 42406
rect 4598 42404 4622 42406
rect 4678 42404 4684 42406
rect 4376 42395 4684 42404
rect 4068 42356 4120 42362
rect 4068 42298 4120 42304
rect 4252 42220 4304 42226
rect 4252 42162 4304 42168
rect 4068 42152 4120 42158
rect 4068 42094 4120 42100
rect 3896 18788 4016 18816
rect 3896 16522 3924 18788
rect 3976 18692 4028 18698
rect 3976 18634 4028 18640
rect 3988 18290 4016 18634
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3792 14544 3844 14550
rect 3712 14504 3792 14532
rect 3792 14486 3844 14492
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 3896 4826 3924 11018
rect 3988 10198 4016 18226
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 4080 2038 4108 42094
rect 4160 41812 4212 41818
rect 4160 41754 4212 41760
rect 4172 41414 4200 41754
rect 4264 41585 4292 42162
rect 4250 41576 4306 41585
rect 4250 41511 4306 41520
rect 4172 41386 4292 41414
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4172 25906 4200 26930
rect 4160 25900 4212 25906
rect 4160 25842 4212 25848
rect 4264 22094 4292 41386
rect 4376 41372 4684 41381
rect 4376 41370 4382 41372
rect 4438 41370 4462 41372
rect 4518 41370 4542 41372
rect 4598 41370 4622 41372
rect 4678 41370 4684 41372
rect 4438 41318 4440 41370
rect 4620 41318 4622 41370
rect 4376 41316 4382 41318
rect 4438 41316 4462 41318
rect 4518 41316 4542 41318
rect 4598 41316 4622 41318
rect 4678 41316 4684 41318
rect 4376 41307 4684 41316
rect 4376 40284 4684 40293
rect 4376 40282 4382 40284
rect 4438 40282 4462 40284
rect 4518 40282 4542 40284
rect 4598 40282 4622 40284
rect 4678 40282 4684 40284
rect 4438 40230 4440 40282
rect 4620 40230 4622 40282
rect 4376 40228 4382 40230
rect 4438 40228 4462 40230
rect 4518 40228 4542 40230
rect 4598 40228 4622 40230
rect 4678 40228 4684 40230
rect 4376 40219 4684 40228
rect 4376 39196 4684 39205
rect 4376 39194 4382 39196
rect 4438 39194 4462 39196
rect 4518 39194 4542 39196
rect 4598 39194 4622 39196
rect 4678 39194 4684 39196
rect 4438 39142 4440 39194
rect 4620 39142 4622 39194
rect 4376 39140 4382 39142
rect 4438 39140 4462 39142
rect 4518 39140 4542 39142
rect 4598 39140 4622 39142
rect 4678 39140 4684 39142
rect 4376 39131 4684 39140
rect 4376 38108 4684 38117
rect 4376 38106 4382 38108
rect 4438 38106 4462 38108
rect 4518 38106 4542 38108
rect 4598 38106 4622 38108
rect 4678 38106 4684 38108
rect 4438 38054 4440 38106
rect 4620 38054 4622 38106
rect 4376 38052 4382 38054
rect 4438 38052 4462 38054
rect 4518 38052 4542 38054
rect 4598 38052 4622 38054
rect 4678 38052 4684 38054
rect 4376 38043 4684 38052
rect 4376 37020 4684 37029
rect 4376 37018 4382 37020
rect 4438 37018 4462 37020
rect 4518 37018 4542 37020
rect 4598 37018 4622 37020
rect 4678 37018 4684 37020
rect 4438 36966 4440 37018
rect 4620 36966 4622 37018
rect 4376 36964 4382 36966
rect 4438 36964 4462 36966
rect 4518 36964 4542 36966
rect 4598 36964 4622 36966
rect 4678 36964 4684 36966
rect 4376 36955 4684 36964
rect 4376 35932 4684 35941
rect 4376 35930 4382 35932
rect 4438 35930 4462 35932
rect 4518 35930 4542 35932
rect 4598 35930 4622 35932
rect 4678 35930 4684 35932
rect 4438 35878 4440 35930
rect 4620 35878 4622 35930
rect 4376 35876 4382 35878
rect 4438 35876 4462 35878
rect 4518 35876 4542 35878
rect 4598 35876 4622 35878
rect 4678 35876 4684 35878
rect 4376 35867 4684 35876
rect 4376 34844 4684 34853
rect 4376 34842 4382 34844
rect 4438 34842 4462 34844
rect 4518 34842 4542 34844
rect 4598 34842 4622 34844
rect 4678 34842 4684 34844
rect 4438 34790 4440 34842
rect 4620 34790 4622 34842
rect 4376 34788 4382 34790
rect 4438 34788 4462 34790
rect 4518 34788 4542 34790
rect 4598 34788 4622 34790
rect 4678 34788 4684 34790
rect 4376 34779 4684 34788
rect 4376 33756 4684 33765
rect 4376 33754 4382 33756
rect 4438 33754 4462 33756
rect 4518 33754 4542 33756
rect 4598 33754 4622 33756
rect 4678 33754 4684 33756
rect 4438 33702 4440 33754
rect 4620 33702 4622 33754
rect 4376 33700 4382 33702
rect 4438 33700 4462 33702
rect 4518 33700 4542 33702
rect 4598 33700 4622 33702
rect 4678 33700 4684 33702
rect 4376 33691 4684 33700
rect 4376 32668 4684 32677
rect 4376 32666 4382 32668
rect 4438 32666 4462 32668
rect 4518 32666 4542 32668
rect 4598 32666 4622 32668
rect 4678 32666 4684 32668
rect 4438 32614 4440 32666
rect 4620 32614 4622 32666
rect 4376 32612 4382 32614
rect 4438 32612 4462 32614
rect 4518 32612 4542 32614
rect 4598 32612 4622 32614
rect 4678 32612 4684 32614
rect 4376 32603 4684 32612
rect 4376 31580 4684 31589
rect 4376 31578 4382 31580
rect 4438 31578 4462 31580
rect 4518 31578 4542 31580
rect 4598 31578 4622 31580
rect 4678 31578 4684 31580
rect 4438 31526 4440 31578
rect 4620 31526 4622 31578
rect 4376 31524 4382 31526
rect 4438 31524 4462 31526
rect 4518 31524 4542 31526
rect 4598 31524 4622 31526
rect 4678 31524 4684 31526
rect 4376 31515 4684 31524
rect 4376 30492 4684 30501
rect 4376 30490 4382 30492
rect 4438 30490 4462 30492
rect 4518 30490 4542 30492
rect 4598 30490 4622 30492
rect 4678 30490 4684 30492
rect 4438 30438 4440 30490
rect 4620 30438 4622 30490
rect 4376 30436 4382 30438
rect 4438 30436 4462 30438
rect 4518 30436 4542 30438
rect 4598 30436 4622 30438
rect 4678 30436 4684 30438
rect 4376 30427 4684 30436
rect 4376 29404 4684 29413
rect 4376 29402 4382 29404
rect 4438 29402 4462 29404
rect 4518 29402 4542 29404
rect 4598 29402 4622 29404
rect 4678 29402 4684 29404
rect 4438 29350 4440 29402
rect 4620 29350 4622 29402
rect 4376 29348 4382 29350
rect 4438 29348 4462 29350
rect 4518 29348 4542 29350
rect 4598 29348 4622 29350
rect 4678 29348 4684 29350
rect 4376 29339 4684 29348
rect 4376 28316 4684 28325
rect 4376 28314 4382 28316
rect 4438 28314 4462 28316
rect 4518 28314 4542 28316
rect 4598 28314 4622 28316
rect 4678 28314 4684 28316
rect 4438 28262 4440 28314
rect 4620 28262 4622 28314
rect 4376 28260 4382 28262
rect 4438 28260 4462 28262
rect 4518 28260 4542 28262
rect 4598 28260 4622 28262
rect 4678 28260 4684 28262
rect 4376 28251 4684 28260
rect 4376 27228 4684 27237
rect 4376 27226 4382 27228
rect 4438 27226 4462 27228
rect 4518 27226 4542 27228
rect 4598 27226 4622 27228
rect 4678 27226 4684 27228
rect 4438 27174 4440 27226
rect 4620 27174 4622 27226
rect 4376 27172 4382 27174
rect 4438 27172 4462 27174
rect 4518 27172 4542 27174
rect 4598 27172 4622 27174
rect 4678 27172 4684 27174
rect 4376 27163 4684 27172
rect 4376 26140 4684 26149
rect 4376 26138 4382 26140
rect 4438 26138 4462 26140
rect 4518 26138 4542 26140
rect 4598 26138 4622 26140
rect 4678 26138 4684 26140
rect 4438 26086 4440 26138
rect 4620 26086 4622 26138
rect 4376 26084 4382 26086
rect 4438 26084 4462 26086
rect 4518 26084 4542 26086
rect 4598 26084 4622 26086
rect 4678 26084 4684 26086
rect 4376 26075 4684 26084
rect 4376 25052 4684 25061
rect 4376 25050 4382 25052
rect 4438 25050 4462 25052
rect 4518 25050 4542 25052
rect 4598 25050 4622 25052
rect 4678 25050 4684 25052
rect 4438 24998 4440 25050
rect 4620 24998 4622 25050
rect 4376 24996 4382 24998
rect 4438 24996 4462 24998
rect 4518 24996 4542 24998
rect 4598 24996 4622 24998
rect 4678 24996 4684 24998
rect 4376 24987 4684 24996
rect 4376 23964 4684 23973
rect 4376 23962 4382 23964
rect 4438 23962 4462 23964
rect 4518 23962 4542 23964
rect 4598 23962 4622 23964
rect 4678 23962 4684 23964
rect 4438 23910 4440 23962
rect 4620 23910 4622 23962
rect 4376 23908 4382 23910
rect 4438 23908 4462 23910
rect 4518 23908 4542 23910
rect 4598 23908 4622 23910
rect 4678 23908 4684 23910
rect 4376 23899 4684 23908
rect 4376 22876 4684 22885
rect 4376 22874 4382 22876
rect 4438 22874 4462 22876
rect 4518 22874 4542 22876
rect 4598 22874 4622 22876
rect 4678 22874 4684 22876
rect 4438 22822 4440 22874
rect 4620 22822 4622 22874
rect 4376 22820 4382 22822
rect 4438 22820 4462 22822
rect 4518 22820 4542 22822
rect 4598 22820 4622 22822
rect 4678 22820 4684 22822
rect 4376 22811 4684 22820
rect 4172 22066 4292 22094
rect 4172 12434 4200 22066
rect 4376 21788 4684 21797
rect 4376 21786 4382 21788
rect 4438 21786 4462 21788
rect 4518 21786 4542 21788
rect 4598 21786 4622 21788
rect 4678 21786 4684 21788
rect 4438 21734 4440 21786
rect 4620 21734 4622 21786
rect 4376 21732 4382 21734
rect 4438 21732 4462 21734
rect 4518 21732 4542 21734
rect 4598 21732 4622 21734
rect 4678 21732 4684 21734
rect 4376 21723 4684 21732
rect 4376 20700 4684 20709
rect 4376 20698 4382 20700
rect 4438 20698 4462 20700
rect 4518 20698 4542 20700
rect 4598 20698 4622 20700
rect 4678 20698 4684 20700
rect 4438 20646 4440 20698
rect 4620 20646 4622 20698
rect 4376 20644 4382 20646
rect 4438 20644 4462 20646
rect 4518 20644 4542 20646
rect 4598 20644 4622 20646
rect 4678 20644 4684 20646
rect 4376 20635 4684 20644
rect 4816 20398 4844 42570
rect 5092 42362 5120 42638
rect 7196 42628 7248 42634
rect 7196 42570 7248 42576
rect 7208 42362 7236 42570
rect 7300 42362 7328 42638
rect 7484 42362 7512 42638
rect 8852 42560 8904 42566
rect 8852 42502 8904 42508
rect 7803 42460 8111 42469
rect 7803 42458 7809 42460
rect 7865 42458 7889 42460
rect 7945 42458 7969 42460
rect 8025 42458 8049 42460
rect 8105 42458 8111 42460
rect 7865 42406 7867 42458
rect 8047 42406 8049 42458
rect 7803 42404 7809 42406
rect 7865 42404 7889 42406
rect 7945 42404 7969 42406
rect 8025 42404 8049 42406
rect 8105 42404 8111 42406
rect 7803 42395 8111 42404
rect 5080 42356 5132 42362
rect 5080 42298 5132 42304
rect 7196 42356 7248 42362
rect 7196 42298 7248 42304
rect 7288 42356 7340 42362
rect 7288 42298 7340 42304
rect 7472 42356 7524 42362
rect 7472 42298 7524 42304
rect 5080 42220 5132 42226
rect 5080 42162 5132 42168
rect 5092 41449 5120 42162
rect 6090 41916 6398 41925
rect 6090 41914 6096 41916
rect 6152 41914 6176 41916
rect 6232 41914 6256 41916
rect 6312 41914 6336 41916
rect 6392 41914 6398 41916
rect 6152 41862 6154 41914
rect 6334 41862 6336 41914
rect 6090 41860 6096 41862
rect 6152 41860 6176 41862
rect 6232 41860 6256 41862
rect 6312 41860 6336 41862
rect 6392 41860 6398 41862
rect 6090 41851 6398 41860
rect 8864 41818 8892 42502
rect 8852 41812 8904 41818
rect 8852 41754 8904 41760
rect 9416 41721 9444 42638
rect 9517 41916 9825 41925
rect 9517 41914 9523 41916
rect 9579 41914 9603 41916
rect 9659 41914 9683 41916
rect 9739 41914 9763 41916
rect 9819 41914 9825 41916
rect 9579 41862 9581 41914
rect 9761 41862 9763 41914
rect 9517 41860 9523 41862
rect 9579 41860 9603 41862
rect 9659 41860 9683 41862
rect 9739 41860 9763 41862
rect 9819 41860 9825 41862
rect 9517 41851 9825 41860
rect 9402 41712 9458 41721
rect 9402 41647 9458 41656
rect 10980 41449 11008 42638
rect 11230 42460 11538 42469
rect 11230 42458 11236 42460
rect 11292 42458 11316 42460
rect 11372 42458 11396 42460
rect 11452 42458 11476 42460
rect 11532 42458 11538 42460
rect 11292 42406 11294 42458
rect 11474 42406 11476 42458
rect 11230 42404 11236 42406
rect 11292 42404 11316 42406
rect 11372 42404 11396 42406
rect 11452 42404 11476 42406
rect 11532 42404 11538 42406
rect 11230 42395 11538 42404
rect 11716 41585 11744 42638
rect 12438 42599 12494 42608
rect 13544 42628 13596 42634
rect 13544 42570 13596 42576
rect 13556 42362 13584 42570
rect 13740 42566 13768 43250
rect 13728 42560 13780 42566
rect 13728 42502 13780 42508
rect 13832 42362 13860 44840
rect 14096 43104 14148 43110
rect 14096 43046 14148 43052
rect 13544 42356 13596 42362
rect 13544 42298 13596 42304
rect 13820 42356 13872 42362
rect 13820 42298 13872 42304
rect 14108 42294 14136 43046
rect 14568 42770 14596 44840
rect 14657 43548 14965 43557
rect 14657 43546 14663 43548
rect 14719 43546 14743 43548
rect 14799 43546 14823 43548
rect 14879 43546 14903 43548
rect 14959 43546 14965 43548
rect 14719 43494 14721 43546
rect 14901 43494 14903 43546
rect 14657 43492 14663 43494
rect 14719 43492 14743 43494
rect 14799 43492 14823 43494
rect 14879 43492 14903 43494
rect 14959 43492 14965 43494
rect 14657 43483 14965 43492
rect 15304 43450 15332 44840
rect 15292 43444 15344 43450
rect 15292 43386 15344 43392
rect 15016 43308 15068 43314
rect 15068 43268 15148 43296
rect 15016 43250 15068 43256
rect 14556 42764 14608 42770
rect 14556 42706 14608 42712
rect 14657 42460 14965 42469
rect 14657 42458 14663 42460
rect 14719 42458 14743 42460
rect 14799 42458 14823 42460
rect 14879 42458 14903 42460
rect 14959 42458 14965 42460
rect 14719 42406 14721 42458
rect 14901 42406 14903 42458
rect 14657 42404 14663 42406
rect 14719 42404 14743 42406
rect 14799 42404 14823 42406
rect 14879 42404 14903 42406
rect 14959 42404 14965 42406
rect 14657 42395 14965 42404
rect 14096 42288 14148 42294
rect 14096 42230 14148 42236
rect 13912 42220 13964 42226
rect 13912 42162 13964 42168
rect 12944 41916 13252 41925
rect 12944 41914 12950 41916
rect 13006 41914 13030 41916
rect 13086 41914 13110 41916
rect 13166 41914 13190 41916
rect 13246 41914 13252 41916
rect 13006 41862 13008 41914
rect 13188 41862 13190 41914
rect 12944 41860 12950 41862
rect 13006 41860 13030 41862
rect 13086 41860 13110 41862
rect 13166 41860 13190 41862
rect 13246 41860 13252 41862
rect 12944 41851 13252 41860
rect 11702 41576 11758 41585
rect 11702 41511 11758 41520
rect 5078 41440 5134 41449
rect 5078 41375 5134 41384
rect 10966 41440 11022 41449
rect 13924 41414 13952 42162
rect 15120 41414 15148 43268
rect 15292 42696 15344 42702
rect 15292 42638 15344 42644
rect 15200 42628 15252 42634
rect 15200 42570 15252 42576
rect 13924 41386 14320 41414
rect 7803 41372 8111 41381
rect 10966 41375 11022 41384
rect 7803 41370 7809 41372
rect 7865 41370 7889 41372
rect 7945 41370 7969 41372
rect 8025 41370 8049 41372
rect 8105 41370 8111 41372
rect 7865 41318 7867 41370
rect 8047 41318 8049 41370
rect 7803 41316 7809 41318
rect 7865 41316 7889 41318
rect 7945 41316 7969 41318
rect 8025 41316 8049 41318
rect 8105 41316 8111 41318
rect 7803 41307 8111 41316
rect 11230 41372 11538 41381
rect 11230 41370 11236 41372
rect 11292 41370 11316 41372
rect 11372 41370 11396 41372
rect 11452 41370 11476 41372
rect 11532 41370 11538 41372
rect 11292 41318 11294 41370
rect 11474 41318 11476 41370
rect 11230 41316 11236 41318
rect 11292 41316 11316 41318
rect 11372 41316 11396 41318
rect 11452 41316 11476 41318
rect 11532 41316 11538 41318
rect 11230 41307 11538 41316
rect 9312 40928 9364 40934
rect 9312 40870 9364 40876
rect 6090 40828 6398 40837
rect 6090 40826 6096 40828
rect 6152 40826 6176 40828
rect 6232 40826 6256 40828
rect 6312 40826 6336 40828
rect 6392 40826 6398 40828
rect 6152 40774 6154 40826
rect 6334 40774 6336 40826
rect 6090 40772 6096 40774
rect 6152 40772 6176 40774
rect 6232 40772 6256 40774
rect 6312 40772 6336 40774
rect 6392 40772 6398 40774
rect 6090 40763 6398 40772
rect 5172 40384 5224 40390
rect 5172 40326 5224 40332
rect 5184 39438 5212 40326
rect 7803 40284 8111 40293
rect 7803 40282 7809 40284
rect 7865 40282 7889 40284
rect 7945 40282 7969 40284
rect 8025 40282 8049 40284
rect 8105 40282 8111 40284
rect 7865 40230 7867 40282
rect 8047 40230 8049 40282
rect 7803 40228 7809 40230
rect 7865 40228 7889 40230
rect 7945 40228 7969 40230
rect 8025 40228 8049 40230
rect 8105 40228 8111 40230
rect 7803 40219 8111 40228
rect 9324 40089 9352 40870
rect 9517 40828 9825 40837
rect 9517 40826 9523 40828
rect 9579 40826 9603 40828
rect 9659 40826 9683 40828
rect 9739 40826 9763 40828
rect 9819 40826 9825 40828
rect 9579 40774 9581 40826
rect 9761 40774 9763 40826
rect 9517 40772 9523 40774
rect 9579 40772 9603 40774
rect 9659 40772 9683 40774
rect 9739 40772 9763 40774
rect 9819 40772 9825 40774
rect 9517 40763 9825 40772
rect 12944 40828 13252 40837
rect 12944 40826 12950 40828
rect 13006 40826 13030 40828
rect 13086 40826 13110 40828
rect 13166 40826 13190 40828
rect 13246 40826 13252 40828
rect 13006 40774 13008 40826
rect 13188 40774 13190 40826
rect 12944 40772 12950 40774
rect 13006 40772 13030 40774
rect 13086 40772 13110 40774
rect 13166 40772 13190 40774
rect 13246 40772 13252 40774
rect 12944 40763 13252 40772
rect 13544 40452 13596 40458
rect 13544 40394 13596 40400
rect 11230 40284 11538 40293
rect 11230 40282 11236 40284
rect 11292 40282 11316 40284
rect 11372 40282 11396 40284
rect 11452 40282 11476 40284
rect 11532 40282 11538 40284
rect 11292 40230 11294 40282
rect 11474 40230 11476 40282
rect 11230 40228 11236 40230
rect 11292 40228 11316 40230
rect 11372 40228 11396 40230
rect 11452 40228 11476 40230
rect 11532 40228 11538 40230
rect 11230 40219 11538 40228
rect 13556 40186 13584 40394
rect 13728 40384 13780 40390
rect 13728 40326 13780 40332
rect 13544 40180 13596 40186
rect 13544 40122 13596 40128
rect 9310 40080 9366 40089
rect 9310 40015 9312 40024
rect 9364 40015 9366 40024
rect 13360 40044 13412 40050
rect 9312 39986 9364 39992
rect 13360 39986 13412 39992
rect 6090 39740 6398 39749
rect 6090 39738 6096 39740
rect 6152 39738 6176 39740
rect 6232 39738 6256 39740
rect 6312 39738 6336 39740
rect 6392 39738 6398 39740
rect 6152 39686 6154 39738
rect 6334 39686 6336 39738
rect 6090 39684 6096 39686
rect 6152 39684 6176 39686
rect 6232 39684 6256 39686
rect 6312 39684 6336 39686
rect 6392 39684 6398 39686
rect 6090 39675 6398 39684
rect 9517 39740 9825 39749
rect 9517 39738 9523 39740
rect 9579 39738 9603 39740
rect 9659 39738 9683 39740
rect 9739 39738 9763 39740
rect 9819 39738 9825 39740
rect 9579 39686 9581 39738
rect 9761 39686 9763 39738
rect 9517 39684 9523 39686
rect 9579 39684 9603 39686
rect 9659 39684 9683 39686
rect 9739 39684 9763 39686
rect 9819 39684 9825 39686
rect 9517 39675 9825 39684
rect 12944 39740 13252 39749
rect 12944 39738 12950 39740
rect 13006 39738 13030 39740
rect 13086 39738 13110 39740
rect 13166 39738 13190 39740
rect 13246 39738 13252 39740
rect 13006 39686 13008 39738
rect 13188 39686 13190 39738
rect 12944 39684 12950 39686
rect 13006 39684 13030 39686
rect 13086 39684 13110 39686
rect 13166 39684 13190 39686
rect 13246 39684 13252 39686
rect 12944 39675 13252 39684
rect 13372 39642 13400 39986
rect 13740 39817 13768 40326
rect 13912 40044 13964 40050
rect 13912 39986 13964 39992
rect 13726 39808 13782 39817
rect 13726 39743 13782 39752
rect 13360 39636 13412 39642
rect 13360 39578 13412 39584
rect 13924 39574 13952 39986
rect 14004 39840 14056 39846
rect 14004 39782 14056 39788
rect 14188 39840 14240 39846
rect 14188 39782 14240 39788
rect 13912 39568 13964 39574
rect 14016 39545 14044 39782
rect 14200 39545 14228 39782
rect 13912 39510 13964 39516
rect 14002 39536 14058 39545
rect 14002 39471 14058 39480
rect 14186 39536 14242 39545
rect 14186 39471 14242 39480
rect 5172 39432 5224 39438
rect 5172 39374 5224 39380
rect 12808 39432 12860 39438
rect 12808 39374 12860 39380
rect 13268 39432 13320 39438
rect 13268 39374 13320 39380
rect 4896 27464 4948 27470
rect 4896 27406 4948 27412
rect 4908 26926 4936 27406
rect 4896 26920 4948 26926
rect 4896 26862 4948 26868
rect 5080 25968 5132 25974
rect 5080 25910 5132 25916
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 4908 23730 4936 24142
rect 4988 24132 5040 24138
rect 4988 24074 5040 24080
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 5000 21690 5028 24074
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4376 19612 4684 19621
rect 4376 19610 4382 19612
rect 4438 19610 4462 19612
rect 4518 19610 4542 19612
rect 4598 19610 4622 19612
rect 4678 19610 4684 19612
rect 4438 19558 4440 19610
rect 4620 19558 4622 19610
rect 4376 19556 4382 19558
rect 4438 19556 4462 19558
rect 4518 19556 4542 19558
rect 4598 19556 4622 19558
rect 4678 19556 4684 19558
rect 4376 19547 4684 19556
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4376 18524 4684 18533
rect 4376 18522 4382 18524
rect 4438 18522 4462 18524
rect 4518 18522 4542 18524
rect 4598 18522 4622 18524
rect 4678 18522 4684 18524
rect 4438 18470 4440 18522
rect 4620 18470 4622 18522
rect 4376 18468 4382 18470
rect 4438 18468 4462 18470
rect 4518 18468 4542 18470
rect 4598 18468 4622 18470
rect 4678 18468 4684 18470
rect 4376 18459 4684 18468
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4264 13870 4292 18158
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 4724 12986 4752 18906
rect 4816 18222 4844 20334
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4172 12406 4752 12434
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4172 9926 4200 10406
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4264 5778 4292 10406
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4724 5574 4752 12406
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4908 11694 4936 12242
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4908 11218 4936 11630
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4908 9042 4936 11154
rect 5000 11082 5028 20538
rect 5092 17218 5120 25910
rect 5184 23730 5212 39374
rect 7803 39196 8111 39205
rect 7803 39194 7809 39196
rect 7865 39194 7889 39196
rect 7945 39194 7969 39196
rect 8025 39194 8049 39196
rect 8105 39194 8111 39196
rect 7865 39142 7867 39194
rect 8047 39142 8049 39194
rect 7803 39140 7809 39142
rect 7865 39140 7889 39142
rect 7945 39140 7969 39142
rect 8025 39140 8049 39142
rect 8105 39140 8111 39142
rect 7803 39131 8111 39140
rect 11230 39196 11538 39205
rect 11230 39194 11236 39196
rect 11292 39194 11316 39196
rect 11372 39194 11396 39196
rect 11452 39194 11476 39196
rect 11532 39194 11538 39196
rect 11292 39142 11294 39194
rect 11474 39142 11476 39194
rect 11230 39140 11236 39142
rect 11292 39140 11316 39142
rect 11372 39140 11396 39142
rect 11452 39140 11476 39142
rect 11532 39140 11538 39142
rect 11230 39131 11538 39140
rect 12820 39030 12848 39374
rect 12808 39024 12860 39030
rect 12808 38966 12860 38972
rect 12716 38956 12768 38962
rect 12716 38898 12768 38904
rect 12348 38888 12400 38894
rect 12348 38830 12400 38836
rect 6090 38652 6398 38661
rect 6090 38650 6096 38652
rect 6152 38650 6176 38652
rect 6232 38650 6256 38652
rect 6312 38650 6336 38652
rect 6392 38650 6398 38652
rect 6152 38598 6154 38650
rect 6334 38598 6336 38650
rect 6090 38596 6096 38598
rect 6152 38596 6176 38598
rect 6232 38596 6256 38598
rect 6312 38596 6336 38598
rect 6392 38596 6398 38598
rect 6090 38587 6398 38596
rect 9517 38652 9825 38661
rect 9517 38650 9523 38652
rect 9579 38650 9603 38652
rect 9659 38650 9683 38652
rect 9739 38650 9763 38652
rect 9819 38650 9825 38652
rect 9579 38598 9581 38650
rect 9761 38598 9763 38650
rect 9517 38596 9523 38598
rect 9579 38596 9603 38598
rect 9659 38596 9683 38598
rect 9739 38596 9763 38598
rect 9819 38596 9825 38598
rect 9517 38587 9825 38596
rect 7803 38108 8111 38117
rect 7803 38106 7809 38108
rect 7865 38106 7889 38108
rect 7945 38106 7969 38108
rect 8025 38106 8049 38108
rect 8105 38106 8111 38108
rect 7865 38054 7867 38106
rect 8047 38054 8049 38106
rect 7803 38052 7809 38054
rect 7865 38052 7889 38054
rect 7945 38052 7969 38054
rect 8025 38052 8049 38054
rect 8105 38052 8111 38054
rect 7803 38043 8111 38052
rect 11230 38108 11538 38117
rect 11230 38106 11236 38108
rect 11292 38106 11316 38108
rect 11372 38106 11396 38108
rect 11452 38106 11476 38108
rect 11532 38106 11538 38108
rect 11292 38054 11294 38106
rect 11474 38054 11476 38106
rect 11230 38052 11236 38054
rect 11292 38052 11316 38054
rect 11372 38052 11396 38054
rect 11452 38052 11476 38054
rect 11532 38052 11538 38054
rect 11230 38043 11538 38052
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 7656 37732 7708 37738
rect 7656 37674 7708 37680
rect 6090 37564 6398 37573
rect 6090 37562 6096 37564
rect 6152 37562 6176 37564
rect 6232 37562 6256 37564
rect 6312 37562 6336 37564
rect 6392 37562 6398 37564
rect 6152 37510 6154 37562
rect 6334 37510 6336 37562
rect 6090 37508 6096 37510
rect 6152 37508 6176 37510
rect 6232 37508 6256 37510
rect 6312 37508 6336 37510
rect 6392 37508 6398 37510
rect 6090 37499 6398 37508
rect 6826 36680 6882 36689
rect 6826 36615 6882 36624
rect 6090 36476 6398 36485
rect 6090 36474 6096 36476
rect 6152 36474 6176 36476
rect 6232 36474 6256 36476
rect 6312 36474 6336 36476
rect 6392 36474 6398 36476
rect 6152 36422 6154 36474
rect 6334 36422 6336 36474
rect 6090 36420 6096 36422
rect 6152 36420 6176 36422
rect 6232 36420 6256 36422
rect 6312 36420 6336 36422
rect 6392 36420 6398 36422
rect 6090 36411 6398 36420
rect 6840 36106 6868 36615
rect 5816 36100 5868 36106
rect 5816 36042 5868 36048
rect 6828 36100 6880 36106
rect 6828 36042 6880 36048
rect 5540 35080 5592 35086
rect 5540 35022 5592 35028
rect 5552 33402 5580 35022
rect 5724 34740 5776 34746
rect 5724 34682 5776 34688
rect 5460 33374 5580 33402
rect 5460 31754 5488 33374
rect 5276 31726 5488 31754
rect 5276 30598 5304 31726
rect 5264 30592 5316 30598
rect 5264 30534 5316 30540
rect 5276 27402 5304 30534
rect 5630 29200 5686 29209
rect 5630 29135 5686 29144
rect 5264 27396 5316 27402
rect 5264 27338 5316 27344
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5184 22234 5212 23666
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5276 17320 5304 27338
rect 5540 24676 5592 24682
rect 5540 24618 5592 24624
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5460 17785 5488 23258
rect 5552 22030 5580 24618
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5644 20754 5672 29135
rect 5552 20726 5672 20754
rect 5552 19990 5580 20726
rect 5736 20618 5764 34682
rect 5828 31754 5856 36042
rect 7196 36032 7248 36038
rect 7196 35974 7248 35980
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 6012 35193 6040 35430
rect 6090 35388 6398 35397
rect 6090 35386 6096 35388
rect 6152 35386 6176 35388
rect 6232 35386 6256 35388
rect 6312 35386 6336 35388
rect 6392 35386 6398 35388
rect 6152 35334 6154 35386
rect 6334 35334 6336 35386
rect 6090 35332 6096 35334
rect 6152 35332 6176 35334
rect 6232 35332 6256 35334
rect 6312 35332 6336 35334
rect 6392 35332 6398 35334
rect 6090 35323 6398 35332
rect 5998 35184 6054 35193
rect 5998 35119 6054 35128
rect 6828 35148 6880 35154
rect 5828 31726 5948 31754
rect 5920 26994 5948 31726
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 6012 24834 6040 35119
rect 6828 35090 6880 35096
rect 6840 34746 6868 35090
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 6828 34740 6880 34746
rect 6828 34682 6880 34688
rect 6090 34300 6398 34309
rect 6090 34298 6096 34300
rect 6152 34298 6176 34300
rect 6232 34298 6256 34300
rect 6312 34298 6336 34300
rect 6392 34298 6398 34300
rect 6152 34246 6154 34298
rect 6334 34246 6336 34298
rect 6090 34244 6096 34246
rect 6152 34244 6176 34246
rect 6232 34244 6256 34246
rect 6312 34244 6336 34246
rect 6392 34244 6398 34246
rect 6090 34235 6398 34244
rect 6090 33212 6398 33221
rect 6090 33210 6096 33212
rect 6152 33210 6176 33212
rect 6232 33210 6256 33212
rect 6312 33210 6336 33212
rect 6392 33210 6398 33212
rect 6152 33158 6154 33210
rect 6334 33158 6336 33210
rect 6090 33156 6096 33158
rect 6152 33156 6176 33158
rect 6232 33156 6256 33158
rect 6312 33156 6336 33158
rect 6392 33156 6398 33158
rect 6090 33147 6398 33156
rect 6460 32768 6512 32774
rect 6460 32710 6512 32716
rect 6090 32124 6398 32133
rect 6090 32122 6096 32124
rect 6152 32122 6176 32124
rect 6232 32122 6256 32124
rect 6312 32122 6336 32124
rect 6392 32122 6398 32124
rect 6152 32070 6154 32122
rect 6334 32070 6336 32122
rect 6090 32068 6096 32070
rect 6152 32068 6176 32070
rect 6232 32068 6256 32070
rect 6312 32068 6336 32070
rect 6392 32068 6398 32070
rect 6090 32059 6398 32068
rect 6472 32026 6500 32710
rect 6932 32450 6960 34954
rect 6932 32434 7052 32450
rect 6920 32428 7052 32434
rect 6972 32422 7052 32428
rect 6920 32370 6972 32376
rect 6918 32328 6974 32337
rect 6918 32263 6974 32272
rect 6460 32020 6512 32026
rect 6460 31962 6512 31968
rect 6472 31754 6500 31962
rect 6644 31884 6696 31890
rect 6644 31826 6696 31832
rect 6472 31726 6592 31754
rect 6564 31686 6592 31726
rect 6552 31680 6604 31686
rect 6552 31622 6604 31628
rect 6656 31414 6684 31826
rect 6932 31754 6960 32263
rect 6920 31748 6972 31754
rect 6920 31690 6972 31696
rect 6644 31408 6696 31414
rect 6644 31350 6696 31356
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 6090 31036 6398 31045
rect 6090 31034 6096 31036
rect 6152 31034 6176 31036
rect 6232 31034 6256 31036
rect 6312 31034 6336 31036
rect 6392 31034 6398 31036
rect 6152 30982 6154 31034
rect 6334 30982 6336 31034
rect 6090 30980 6096 30982
rect 6152 30980 6176 30982
rect 6232 30980 6256 30982
rect 6312 30980 6336 30982
rect 6392 30980 6398 30982
rect 6090 30971 6398 30980
rect 6736 30932 6788 30938
rect 6736 30874 6788 30880
rect 6644 30388 6696 30394
rect 6644 30330 6696 30336
rect 6552 30252 6604 30258
rect 6552 30194 6604 30200
rect 6090 29948 6398 29957
rect 6090 29946 6096 29948
rect 6152 29946 6176 29948
rect 6232 29946 6256 29948
rect 6312 29946 6336 29948
rect 6392 29946 6398 29948
rect 6152 29894 6154 29946
rect 6334 29894 6336 29946
rect 6090 29892 6096 29894
rect 6152 29892 6176 29894
rect 6232 29892 6256 29894
rect 6312 29892 6336 29894
rect 6392 29892 6398 29894
rect 6090 29883 6398 29892
rect 6090 28860 6398 28869
rect 6090 28858 6096 28860
rect 6152 28858 6176 28860
rect 6232 28858 6256 28860
rect 6312 28858 6336 28860
rect 6392 28858 6398 28860
rect 6152 28806 6154 28858
rect 6334 28806 6336 28858
rect 6090 28804 6096 28806
rect 6152 28804 6176 28806
rect 6232 28804 6256 28806
rect 6312 28804 6336 28806
rect 6392 28804 6398 28806
rect 6090 28795 6398 28804
rect 6090 27772 6398 27781
rect 6090 27770 6096 27772
rect 6152 27770 6176 27772
rect 6232 27770 6256 27772
rect 6312 27770 6336 27772
rect 6392 27770 6398 27772
rect 6152 27718 6154 27770
rect 6334 27718 6336 27770
rect 6090 27716 6096 27718
rect 6152 27716 6176 27718
rect 6232 27716 6256 27718
rect 6312 27716 6336 27718
rect 6392 27716 6398 27718
rect 6090 27707 6398 27716
rect 6460 26988 6512 26994
rect 6460 26930 6512 26936
rect 6090 26684 6398 26693
rect 6090 26682 6096 26684
rect 6152 26682 6176 26684
rect 6232 26682 6256 26684
rect 6312 26682 6336 26684
rect 6392 26682 6398 26684
rect 6152 26630 6154 26682
rect 6334 26630 6336 26682
rect 6090 26628 6096 26630
rect 6152 26628 6176 26630
rect 6232 26628 6256 26630
rect 6312 26628 6336 26630
rect 6392 26628 6398 26630
rect 6090 26619 6398 26628
rect 6090 25596 6398 25605
rect 6090 25594 6096 25596
rect 6152 25594 6176 25596
rect 6232 25594 6256 25596
rect 6312 25594 6336 25596
rect 6392 25594 6398 25596
rect 6152 25542 6154 25594
rect 6334 25542 6336 25594
rect 6090 25540 6096 25542
rect 6152 25540 6176 25542
rect 6232 25540 6256 25542
rect 6312 25540 6336 25542
rect 6392 25540 6398 25542
rect 6090 25531 6398 25540
rect 5644 20590 5764 20618
rect 5828 24806 6040 24834
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5552 19417 5580 19926
rect 5538 19408 5594 19417
rect 5538 19343 5594 19352
rect 5644 18766 5672 20590
rect 5828 19990 5856 24806
rect 5908 24744 5960 24750
rect 5908 24686 5960 24692
rect 5920 24313 5948 24686
rect 6090 24508 6398 24517
rect 6090 24506 6096 24508
rect 6152 24506 6176 24508
rect 6232 24506 6256 24508
rect 6312 24506 6336 24508
rect 6392 24506 6398 24508
rect 6152 24454 6154 24506
rect 6334 24454 6336 24506
rect 6090 24452 6096 24454
rect 6152 24452 6176 24454
rect 6232 24452 6256 24454
rect 6312 24452 6336 24454
rect 6392 24452 6398 24454
rect 6090 24443 6398 24452
rect 5906 24304 5962 24313
rect 5906 24239 5962 24248
rect 5920 22030 5948 24239
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 6380 23662 6408 24142
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 5920 21486 5948 21966
rect 5908 21480 5960 21486
rect 5908 21422 5960 21428
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5446 17776 5502 17785
rect 5446 17711 5502 17720
rect 5276 17292 5488 17320
rect 5092 17190 5304 17218
rect 5170 17096 5226 17105
rect 5170 17031 5226 17040
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5092 14482 5120 15438
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5184 11830 5212 17031
rect 5276 11898 5304 17190
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5368 15366 5396 15642
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5460 13802 5488 17292
rect 5736 16640 5764 19110
rect 5828 18698 5856 19790
rect 5816 18692 5868 18698
rect 5816 18634 5868 18640
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5828 17814 5856 18158
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5736 16612 5856 16640
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5552 13394 5580 14418
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4908 7954 4936 8978
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8401 5488 8774
rect 5446 8392 5502 8401
rect 5446 8327 5502 8336
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 5644 7546 5672 14486
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 5736 2774 5764 16458
rect 5828 13938 5856 16612
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5828 13326 5856 13738
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5828 6322 5856 13262
rect 5920 12306 5948 21422
rect 6012 19174 6040 23598
rect 6090 23420 6398 23429
rect 6090 23418 6096 23420
rect 6152 23418 6176 23420
rect 6232 23418 6256 23420
rect 6312 23418 6336 23420
rect 6392 23418 6398 23420
rect 6152 23366 6154 23418
rect 6334 23366 6336 23418
rect 6090 23364 6096 23366
rect 6152 23364 6176 23366
rect 6232 23364 6256 23366
rect 6312 23364 6336 23366
rect 6392 23364 6398 23366
rect 6090 23355 6398 23364
rect 6090 22332 6398 22341
rect 6090 22330 6096 22332
rect 6152 22330 6176 22332
rect 6232 22330 6256 22332
rect 6312 22330 6336 22332
rect 6392 22330 6398 22332
rect 6152 22278 6154 22330
rect 6334 22278 6336 22330
rect 6090 22276 6096 22278
rect 6152 22276 6176 22278
rect 6232 22276 6256 22278
rect 6312 22276 6336 22278
rect 6392 22276 6398 22278
rect 6090 22267 6398 22276
rect 6472 22094 6500 26930
rect 6564 24886 6592 30194
rect 6656 28558 6684 30330
rect 6644 28552 6696 28558
rect 6644 28494 6696 28500
rect 6748 27418 6776 30874
rect 6840 28762 6868 31282
rect 7024 30802 7052 32422
rect 7208 31890 7236 35974
rect 7288 32768 7340 32774
rect 7288 32710 7340 32716
rect 7300 32434 7328 32710
rect 7288 32428 7340 32434
rect 7288 32370 7340 32376
rect 7196 31884 7248 31890
rect 7196 31826 7248 31832
rect 7300 31754 7328 32370
rect 7472 31816 7524 31822
rect 7472 31758 7524 31764
rect 7196 31748 7248 31754
rect 7300 31726 7420 31754
rect 7196 31690 7248 31696
rect 7012 30796 7064 30802
rect 7012 30738 7064 30744
rect 7012 30252 7064 30258
rect 6932 30212 7012 30240
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 6840 28082 6868 28698
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6656 27390 6776 27418
rect 6552 24880 6604 24886
rect 6552 24822 6604 24828
rect 6656 24818 6684 27390
rect 6840 27334 6868 27474
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6748 26926 6776 27270
rect 6840 26926 6868 27270
rect 6736 26920 6788 26926
rect 6736 26862 6788 26868
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6472 22066 6592 22094
rect 6276 22024 6328 22030
rect 6276 21966 6328 21972
rect 6288 21593 6316 21966
rect 6274 21584 6330 21593
rect 6274 21519 6330 21528
rect 6090 21244 6398 21253
rect 6090 21242 6096 21244
rect 6152 21242 6176 21244
rect 6232 21242 6256 21244
rect 6312 21242 6336 21244
rect 6392 21242 6398 21244
rect 6152 21190 6154 21242
rect 6334 21190 6336 21242
rect 6090 21188 6096 21190
rect 6152 21188 6176 21190
rect 6232 21188 6256 21190
rect 6312 21188 6336 21190
rect 6392 21188 6398 21190
rect 6090 21179 6398 21188
rect 6564 21078 6592 22066
rect 6552 21072 6604 21078
rect 6552 21014 6604 21020
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6090 20156 6398 20165
rect 6090 20154 6096 20156
rect 6152 20154 6176 20156
rect 6232 20154 6256 20156
rect 6312 20154 6336 20156
rect 6392 20154 6398 20156
rect 6152 20102 6154 20154
rect 6334 20102 6336 20154
rect 6090 20100 6096 20102
rect 6152 20100 6176 20102
rect 6232 20100 6256 20102
rect 6312 20100 6336 20102
rect 6392 20100 6398 20102
rect 6090 20091 6398 20100
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6090 19068 6398 19077
rect 6090 19066 6096 19068
rect 6152 19066 6176 19068
rect 6232 19066 6256 19068
rect 6312 19066 6336 19068
rect 6392 19066 6398 19068
rect 6152 19014 6154 19066
rect 6334 19014 6336 19066
rect 6090 19012 6096 19014
rect 6152 19012 6176 19014
rect 6232 19012 6256 19014
rect 6312 19012 6336 19014
rect 6392 19012 6398 19014
rect 6090 19003 6398 19012
rect 6000 18692 6052 18698
rect 6000 18634 6052 18640
rect 6012 18086 6040 18634
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 6012 17678 6040 18022
rect 6090 17980 6398 17989
rect 6090 17978 6096 17980
rect 6152 17978 6176 17980
rect 6232 17978 6256 17980
rect 6312 17978 6336 17980
rect 6392 17978 6398 17980
rect 6152 17926 6154 17978
rect 6334 17926 6336 17978
rect 6090 17924 6096 17926
rect 6152 17924 6176 17926
rect 6232 17924 6256 17926
rect 6312 17924 6336 17926
rect 6392 17924 6398 17926
rect 6090 17915 6398 17924
rect 6472 17728 6500 20878
rect 6564 17898 6592 20878
rect 6656 18222 6684 24754
rect 6748 24342 6776 26862
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 6736 24200 6788 24206
rect 6736 24142 6788 24148
rect 6748 23746 6776 24142
rect 6840 23866 6868 26862
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6748 23718 6868 23746
rect 6840 21622 6868 23718
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6736 21072 6788 21078
rect 6736 21014 6788 21020
rect 6748 20806 6776 21014
rect 6932 21010 6960 30212
rect 7012 30194 7064 30200
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6932 19854 6960 20946
rect 7024 20913 7052 29038
rect 7104 27872 7156 27878
rect 7104 27814 7156 27820
rect 7116 26790 7144 27814
rect 7104 26784 7156 26790
rect 7104 26726 7156 26732
rect 7116 26586 7144 26726
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 7116 24206 7144 25230
rect 7208 24954 7236 31690
rect 7288 30592 7340 30598
rect 7288 30534 7340 30540
rect 7300 30054 7328 30534
rect 7288 30048 7340 30054
rect 7288 29990 7340 29996
rect 7288 29028 7340 29034
rect 7288 28970 7340 28976
rect 7300 27674 7328 28970
rect 7392 28762 7420 31726
rect 7484 30326 7512 31758
rect 7564 31408 7616 31414
rect 7564 31350 7616 31356
rect 7472 30320 7524 30326
rect 7472 30262 7524 30268
rect 7380 28756 7432 28762
rect 7380 28698 7432 28704
rect 7392 28218 7420 28698
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 7380 28212 7432 28218
rect 7380 28154 7432 28160
rect 7288 27668 7340 27674
rect 7288 27610 7340 27616
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7116 23905 7144 24142
rect 7194 24032 7250 24041
rect 7194 23967 7250 23976
rect 7102 23896 7158 23905
rect 7102 23831 7158 23840
rect 7208 23322 7236 23967
rect 7300 23730 7328 27610
rect 7484 27470 7512 28358
rect 7576 28150 7604 31350
rect 7564 28144 7616 28150
rect 7564 28086 7616 28092
rect 7668 27614 7696 37674
rect 9517 37564 9825 37573
rect 9517 37562 9523 37564
rect 9579 37562 9603 37564
rect 9659 37562 9683 37564
rect 9739 37562 9763 37564
rect 9819 37562 9825 37564
rect 9579 37510 9581 37562
rect 9761 37510 9763 37562
rect 9517 37508 9523 37510
rect 9579 37508 9603 37510
rect 9659 37508 9683 37510
rect 9739 37508 9763 37510
rect 9819 37508 9825 37510
rect 9517 37499 9825 37508
rect 10796 37466 10824 37810
rect 12256 37732 12308 37738
rect 12256 37674 12308 37680
rect 10784 37460 10836 37466
rect 10784 37402 10836 37408
rect 10508 37324 10560 37330
rect 10508 37266 10560 37272
rect 9862 37224 9918 37233
rect 9128 37188 9180 37194
rect 9862 37159 9918 37168
rect 9128 37130 9180 37136
rect 7803 37020 8111 37029
rect 7803 37018 7809 37020
rect 7865 37018 7889 37020
rect 7945 37018 7969 37020
rect 8025 37018 8049 37020
rect 8105 37018 8111 37020
rect 7865 36966 7867 37018
rect 8047 36966 8049 37018
rect 7803 36964 7809 36966
rect 7865 36964 7889 36966
rect 7945 36964 7969 36966
rect 8025 36964 8049 36966
rect 8105 36964 8111 36966
rect 7803 36955 8111 36964
rect 9140 36378 9168 37130
rect 9517 36476 9825 36485
rect 9517 36474 9523 36476
rect 9579 36474 9603 36476
rect 9659 36474 9683 36476
rect 9739 36474 9763 36476
rect 9819 36474 9825 36476
rect 9579 36422 9581 36474
rect 9761 36422 9763 36474
rect 9517 36420 9523 36422
rect 9579 36420 9603 36422
rect 9659 36420 9683 36422
rect 9739 36420 9763 36422
rect 9819 36420 9825 36422
rect 9517 36411 9825 36420
rect 9128 36372 9180 36378
rect 9128 36314 9180 36320
rect 9312 36168 9364 36174
rect 9312 36110 9364 36116
rect 8300 36100 8352 36106
rect 8300 36042 8352 36048
rect 7803 35932 8111 35941
rect 7803 35930 7809 35932
rect 7865 35930 7889 35932
rect 7945 35930 7969 35932
rect 8025 35930 8049 35932
rect 8105 35930 8111 35932
rect 7865 35878 7867 35930
rect 8047 35878 8049 35930
rect 7803 35876 7809 35878
rect 7865 35876 7889 35878
rect 7945 35876 7969 35878
rect 8025 35876 8049 35878
rect 8105 35876 8111 35878
rect 7803 35867 8111 35876
rect 7803 34844 8111 34853
rect 7803 34842 7809 34844
rect 7865 34842 7889 34844
rect 7945 34842 7969 34844
rect 8025 34842 8049 34844
rect 8105 34842 8111 34844
rect 7865 34790 7867 34842
rect 8047 34790 8049 34842
rect 7803 34788 7809 34790
rect 7865 34788 7889 34790
rect 7945 34788 7969 34790
rect 8025 34788 8049 34790
rect 8105 34788 8111 34790
rect 7803 34779 8111 34788
rect 7803 33756 8111 33765
rect 7803 33754 7809 33756
rect 7865 33754 7889 33756
rect 7945 33754 7969 33756
rect 8025 33754 8049 33756
rect 8105 33754 8111 33756
rect 7865 33702 7867 33754
rect 8047 33702 8049 33754
rect 7803 33700 7809 33702
rect 7865 33700 7889 33702
rect 7945 33700 7969 33702
rect 8025 33700 8049 33702
rect 8105 33700 8111 33702
rect 7803 33691 8111 33700
rect 7803 32668 8111 32677
rect 7803 32666 7809 32668
rect 7865 32666 7889 32668
rect 7945 32666 7969 32668
rect 8025 32666 8049 32668
rect 8105 32666 8111 32668
rect 7865 32614 7867 32666
rect 8047 32614 8049 32666
rect 7803 32612 7809 32614
rect 7865 32612 7889 32614
rect 7945 32612 7969 32614
rect 8025 32612 8049 32614
rect 8105 32612 8111 32614
rect 7803 32603 8111 32612
rect 8024 32224 8076 32230
rect 8024 32166 8076 32172
rect 8036 31754 8064 32166
rect 8312 32026 8340 36042
rect 9324 35834 9352 36110
rect 9312 35828 9364 35834
rect 9312 35770 9364 35776
rect 8576 35692 8628 35698
rect 8576 35634 8628 35640
rect 8484 32836 8536 32842
rect 8484 32778 8536 32784
rect 8496 32502 8524 32778
rect 8484 32496 8536 32502
rect 8484 32438 8536 32444
rect 8300 32020 8352 32026
rect 8300 31962 8352 31968
rect 8496 31754 8524 32438
rect 8036 31726 8248 31754
rect 7803 31580 8111 31589
rect 7803 31578 7809 31580
rect 7865 31578 7889 31580
rect 7945 31578 7969 31580
rect 8025 31578 8049 31580
rect 8105 31578 8111 31580
rect 7865 31526 7867 31578
rect 8047 31526 8049 31578
rect 7803 31524 7809 31526
rect 7865 31524 7889 31526
rect 7945 31524 7969 31526
rect 8025 31524 8049 31526
rect 8105 31524 8111 31526
rect 7803 31515 8111 31524
rect 7803 30492 8111 30501
rect 7803 30490 7809 30492
rect 7865 30490 7889 30492
rect 7945 30490 7969 30492
rect 8025 30490 8049 30492
rect 8105 30490 8111 30492
rect 7865 30438 7867 30490
rect 8047 30438 8049 30490
rect 7803 30436 7809 30438
rect 7865 30436 7889 30438
rect 7945 30436 7969 30438
rect 8025 30436 8049 30438
rect 8105 30436 8111 30438
rect 7803 30427 8111 30436
rect 8116 30184 8168 30190
rect 8116 30126 8168 30132
rect 8128 29850 8156 30126
rect 8116 29844 8168 29850
rect 8116 29786 8168 29792
rect 7803 29404 8111 29413
rect 7803 29402 7809 29404
rect 7865 29402 7889 29404
rect 7945 29402 7969 29404
rect 8025 29402 8049 29404
rect 8105 29402 8111 29404
rect 7865 29350 7867 29402
rect 8047 29350 8049 29402
rect 7803 29348 7809 29350
rect 7865 29348 7889 29350
rect 7945 29348 7969 29350
rect 8025 29348 8049 29350
rect 8105 29348 8111 29350
rect 7803 29339 8111 29348
rect 8220 29345 8248 31726
rect 8312 31726 8524 31754
rect 8206 29336 8262 29345
rect 8206 29271 8262 29280
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 7803 28316 8111 28325
rect 7803 28314 7809 28316
rect 7865 28314 7889 28316
rect 7945 28314 7969 28316
rect 8025 28314 8049 28316
rect 8105 28314 8111 28316
rect 7865 28262 7867 28314
rect 8047 28262 8049 28314
rect 7803 28260 7809 28262
rect 7865 28260 7889 28262
rect 7945 28260 7969 28262
rect 8025 28260 8049 28262
rect 8105 28260 8111 28262
rect 7803 28251 8111 28260
rect 8116 27872 8168 27878
rect 8116 27814 8168 27820
rect 7576 27586 7696 27614
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 7472 26444 7524 26450
rect 7392 26404 7472 26432
rect 7392 25294 7420 26404
rect 7472 26386 7524 26392
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7392 24818 7420 25230
rect 7576 24818 7604 27586
rect 8128 27538 8156 27814
rect 7840 27532 7892 27538
rect 7840 27474 7892 27480
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 7852 27316 7880 27474
rect 8220 27334 8248 28902
rect 7742 27288 7880 27316
rect 8208 27328 8260 27334
rect 7742 27112 7770 27288
rect 8208 27270 8260 27276
rect 7803 27228 8111 27237
rect 7803 27226 7809 27228
rect 7865 27226 7889 27228
rect 7945 27226 7969 27228
rect 8025 27226 8049 27228
rect 8105 27226 8111 27228
rect 7865 27174 7867 27226
rect 8047 27174 8049 27226
rect 7803 27172 7809 27174
rect 7865 27172 7889 27174
rect 7945 27172 7969 27174
rect 8025 27172 8049 27174
rect 8105 27172 8111 27174
rect 7803 27163 8111 27172
rect 7742 27084 7788 27112
rect 7760 26926 7788 27084
rect 7748 26920 7800 26926
rect 7668 26880 7748 26908
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7380 24676 7432 24682
rect 7380 24618 7432 24624
rect 7392 24410 7420 24618
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7484 24410 7512 24550
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7668 24290 7696 26880
rect 7748 26862 7800 26868
rect 7932 26920 7984 26926
rect 7932 26862 7984 26868
rect 7944 26586 7972 26862
rect 7932 26580 7984 26586
rect 7932 26522 7984 26528
rect 7803 26140 8111 26149
rect 7803 26138 7809 26140
rect 7865 26138 7889 26140
rect 7945 26138 7969 26140
rect 8025 26138 8049 26140
rect 8105 26138 8111 26140
rect 7865 26086 7867 26138
rect 8047 26086 8049 26138
rect 7803 26084 7809 26086
rect 7865 26084 7889 26086
rect 7945 26084 7969 26086
rect 8025 26084 8049 26086
rect 8105 26084 8111 26086
rect 7803 26075 8111 26084
rect 8208 25288 8260 25294
rect 8206 25256 8208 25265
rect 8260 25256 8262 25265
rect 8206 25191 8262 25200
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 7803 25052 8111 25061
rect 7803 25050 7809 25052
rect 7865 25050 7889 25052
rect 7945 25050 7969 25052
rect 8025 25050 8049 25052
rect 8105 25050 8111 25052
rect 7865 24998 7867 25050
rect 8047 24998 8049 25050
rect 7803 24996 7809 24998
rect 7865 24996 7889 24998
rect 7945 24996 7969 24998
rect 8025 24996 8049 24998
rect 8105 24996 8111 24998
rect 7803 24987 8111 24996
rect 7748 24948 7800 24954
rect 7748 24890 7800 24896
rect 7392 24262 7696 24290
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7300 23322 7328 23666
rect 7392 23662 7420 24262
rect 7760 24154 7788 24890
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7852 24206 7880 24550
rect 7668 24126 7788 24154
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7576 23730 7604 24006
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7392 23202 7420 23598
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7300 23174 7420 23202
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7010 20904 7066 20913
rect 7010 20839 7066 20848
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6748 18714 6776 19382
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6840 18884 6868 19314
rect 6920 18896 6972 18902
rect 6840 18856 6920 18884
rect 6920 18838 6972 18844
rect 6748 18686 6868 18714
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 18306 6776 18566
rect 6840 18426 6868 18686
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6748 18278 6868 18306
rect 6644 18216 6696 18222
rect 6696 18176 6776 18204
rect 6644 18158 6696 18164
rect 6564 17870 6684 17898
rect 6472 17700 6592 17728
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6458 17640 6514 17649
rect 6012 16658 6040 17614
rect 6458 17575 6460 17584
rect 6512 17575 6514 17584
rect 6460 17546 6512 17552
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6564 16454 6592 17700
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6380 15094 6408 15574
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6368 15088 6420 15094
rect 6368 15030 6420 15036
rect 6472 14958 6500 15302
rect 6564 15162 6592 16390
rect 6656 16250 6684 17870
rect 6748 16794 6776 18176
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 6656 12170 6684 16050
rect 6748 16046 6776 16594
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6748 11098 6776 15098
rect 6840 12850 6868 18278
rect 7024 17954 7052 20198
rect 7116 19938 7144 21558
rect 7300 20924 7328 23174
rect 7484 21622 7512 23258
rect 7564 22024 7616 22030
rect 7562 21992 7564 22001
rect 7616 21992 7618 22001
rect 7562 21927 7618 21936
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7392 21146 7420 21286
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7380 20936 7432 20942
rect 7208 20896 7380 20924
rect 7208 20262 7236 20896
rect 7380 20878 7432 20884
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7300 19990 7328 20402
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7288 19984 7340 19990
rect 7116 19910 7236 19938
rect 7288 19926 7340 19932
rect 7104 19848 7156 19854
rect 7208 19836 7236 19910
rect 7208 19808 7328 19836
rect 7104 19790 7156 19796
rect 7116 19514 7144 19790
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 19514 7236 19654
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7196 19315 7248 19321
rect 7196 19257 7248 19263
rect 7208 18902 7236 19257
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 6932 17926 7052 17954
rect 6932 15978 6960 17926
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 7024 17202 7052 17818
rect 7116 17678 7144 18566
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17338 7236 17478
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7300 17218 7328 19808
rect 7392 19310 7420 20198
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7378 18864 7434 18873
rect 7378 18799 7434 18808
rect 7392 18766 7420 18799
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7208 17190 7328 17218
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6932 15638 6960 15914
rect 6920 15632 6972 15638
rect 6920 15574 6972 15580
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6932 14618 6960 14962
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7024 14362 7052 17138
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7116 16454 7144 16730
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7116 15026 7144 16186
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7208 14550 7236 17190
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7102 14376 7158 14385
rect 7024 14334 7102 14362
rect 7102 14311 7158 14320
rect 7104 14272 7156 14278
rect 7024 14232 7104 14260
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 7024 12434 7052 14232
rect 7104 14214 7156 14220
rect 7104 14068 7156 14074
rect 7208 14056 7236 14486
rect 7156 14028 7236 14056
rect 7104 14010 7156 14016
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7102 13696 7158 13705
rect 7102 13631 7158 13640
rect 7116 12918 7144 13631
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7024 12406 7144 12434
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 11218 6868 11630
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10606 6500 10950
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 6472 10062 6500 10542
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6564 9654 6592 11086
rect 6748 11070 6868 11098
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6656 10674 6684 10950
rect 6748 10742 6776 10950
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6840 10606 6868 11070
rect 6828 10600 6880 10606
rect 6826 10568 6828 10577
rect 6880 10568 6882 10577
rect 6932 10538 6960 11494
rect 7024 10810 7052 11494
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7116 10690 7144 12406
rect 7024 10662 7144 10690
rect 6826 10503 6882 10512
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 10266 6868 10406
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 6472 9178 6500 9522
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6564 9178 6592 9318
rect 6656 9178 6684 9930
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6656 8634 6684 8910
rect 6932 8634 6960 9522
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 5736 2746 5856 2774
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 5828 2106 5856 2746
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 6564 2106 6592 7482
rect 6932 7342 6960 7754
rect 7024 7410 7052 10662
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7116 8974 7144 9522
rect 7104 8968 7156 8974
rect 7102 8936 7104 8945
rect 7156 8936 7158 8945
rect 7102 8871 7158 8880
rect 7208 8537 7236 13806
rect 7300 11694 7328 17070
rect 7392 13734 7420 18702
rect 7484 18290 7512 21558
rect 7576 20942 7604 21830
rect 7668 21146 7696 24126
rect 7944 24052 7972 24686
rect 7742 24024 7972 24052
rect 7742 23848 7770 24024
rect 7803 23964 8111 23973
rect 7803 23962 7809 23964
rect 7865 23962 7889 23964
rect 7945 23962 7969 23964
rect 8025 23962 8049 23964
rect 8105 23962 8111 23964
rect 7865 23910 7867 23962
rect 8047 23910 8049 23962
rect 7803 23908 7809 23910
rect 7865 23908 7889 23910
rect 7945 23908 7969 23910
rect 8025 23908 8049 23910
rect 8105 23908 8111 23910
rect 7803 23899 8111 23908
rect 8220 23866 8248 25094
rect 8208 23860 8260 23866
rect 7742 23820 7788 23848
rect 7760 23032 7788 23820
rect 8208 23802 8260 23808
rect 7742 23004 7788 23032
rect 7742 22760 7770 23004
rect 7803 22876 8111 22885
rect 7803 22874 7809 22876
rect 7865 22874 7889 22876
rect 7945 22874 7969 22876
rect 8025 22874 8049 22876
rect 8105 22874 8111 22876
rect 7865 22822 7867 22874
rect 8047 22822 8049 22874
rect 7803 22820 7809 22822
rect 7865 22820 7889 22822
rect 7945 22820 7969 22822
rect 8025 22820 8049 22822
rect 8105 22820 8111 22822
rect 7803 22811 8111 22820
rect 7742 22732 7788 22760
rect 7760 22574 7788 22732
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7760 22234 7788 22510
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7760 21876 7788 22170
rect 7742 21848 7788 21876
rect 7742 21672 7770 21848
rect 7803 21788 8111 21797
rect 7803 21786 7809 21788
rect 7865 21786 7889 21788
rect 7945 21786 7969 21788
rect 8025 21786 8049 21788
rect 8105 21786 8111 21788
rect 7865 21734 7867 21786
rect 8047 21734 8049 21786
rect 7803 21732 7809 21734
rect 7865 21732 7889 21734
rect 7945 21732 7969 21734
rect 8025 21732 8049 21734
rect 8105 21732 8111 21734
rect 7803 21723 8111 21732
rect 7742 21644 7788 21672
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7760 21026 7788 21644
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 7668 20998 7788 21026
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7668 20856 7696 20998
rect 7650 20828 7696 20856
rect 7650 20788 7678 20828
rect 7852 20788 7880 21422
rect 7944 21010 7972 21558
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8036 21078 8064 21422
rect 8208 21344 8260 21350
rect 8312 21332 8340 31726
rect 8484 31340 8536 31346
rect 8484 31282 8536 31288
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8404 29102 8432 30534
rect 8496 30274 8524 31282
rect 8588 30394 8616 35634
rect 9517 35388 9825 35397
rect 9517 35386 9523 35388
rect 9579 35386 9603 35388
rect 9659 35386 9683 35388
rect 9739 35386 9763 35388
rect 9819 35386 9825 35388
rect 9579 35334 9581 35386
rect 9761 35334 9763 35386
rect 9517 35332 9523 35334
rect 9579 35332 9603 35334
rect 9659 35332 9683 35334
rect 9739 35332 9763 35334
rect 9819 35332 9825 35334
rect 9517 35323 9825 35332
rect 9517 34300 9825 34309
rect 9517 34298 9523 34300
rect 9579 34298 9603 34300
rect 9659 34298 9683 34300
rect 9739 34298 9763 34300
rect 9819 34298 9825 34300
rect 9579 34246 9581 34298
rect 9761 34246 9763 34298
rect 9517 34244 9523 34246
rect 9579 34244 9603 34246
rect 9659 34244 9683 34246
rect 9739 34244 9763 34246
rect 9819 34244 9825 34246
rect 9517 34235 9825 34244
rect 8760 33992 8812 33998
rect 8760 33934 8812 33940
rect 8668 32564 8720 32570
rect 8668 32506 8720 32512
rect 8680 30802 8708 32506
rect 8668 30796 8720 30802
rect 8668 30738 8720 30744
rect 8772 30682 8800 33934
rect 9876 33862 9904 37159
rect 10140 36712 10192 36718
rect 10140 36654 10192 36660
rect 10046 36272 10102 36281
rect 10046 36207 10102 36216
rect 9864 33856 9916 33862
rect 9864 33798 9916 33804
rect 9517 33212 9825 33221
rect 9517 33210 9523 33212
rect 9579 33210 9603 33212
rect 9659 33210 9683 33212
rect 9739 33210 9763 33212
rect 9819 33210 9825 33212
rect 9579 33158 9581 33210
rect 9761 33158 9763 33210
rect 9517 33156 9523 33158
rect 9579 33156 9603 33158
rect 9659 33156 9683 33158
rect 9739 33156 9763 33158
rect 9819 33156 9825 33158
rect 9517 33147 9825 33156
rect 10060 33114 10088 36207
rect 10152 35834 10180 36654
rect 10520 36009 10548 37266
rect 11230 37020 11538 37029
rect 11230 37018 11236 37020
rect 11292 37018 11316 37020
rect 11372 37018 11396 37020
rect 11452 37018 11476 37020
rect 11532 37018 11538 37020
rect 11292 36966 11294 37018
rect 11474 36966 11476 37018
rect 11230 36964 11236 36966
rect 11292 36964 11316 36966
rect 11372 36964 11396 36966
rect 11452 36964 11476 36966
rect 11532 36964 11538 36966
rect 11230 36955 11538 36964
rect 11060 36780 11112 36786
rect 11060 36722 11112 36728
rect 12164 36780 12216 36786
rect 12164 36722 12216 36728
rect 10966 36136 11022 36145
rect 10888 36094 10966 36122
rect 10506 36000 10562 36009
rect 10506 35935 10562 35944
rect 10140 35828 10192 35834
rect 10140 35770 10192 35776
rect 10232 35760 10284 35766
rect 10232 35702 10284 35708
rect 10244 34202 10272 35702
rect 10324 35692 10376 35698
rect 10324 35634 10376 35640
rect 10336 35290 10364 35634
rect 10324 35284 10376 35290
rect 10324 35226 10376 35232
rect 10506 35048 10562 35057
rect 10506 34983 10562 34992
rect 10416 34944 10468 34950
rect 10416 34886 10468 34892
rect 10428 34746 10456 34886
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10520 34626 10548 34983
rect 10428 34598 10548 34626
rect 10690 34640 10746 34649
rect 10600 34604 10652 34610
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 10324 33856 10376 33862
rect 10324 33798 10376 33804
rect 10140 33312 10192 33318
rect 10140 33254 10192 33260
rect 10048 33108 10100 33114
rect 10048 33050 10100 33056
rect 8944 32904 8996 32910
rect 8944 32846 8996 32852
rect 8956 32026 8984 32846
rect 9864 32564 9916 32570
rect 9864 32506 9916 32512
rect 9404 32224 9456 32230
rect 9404 32166 9456 32172
rect 8944 32020 8996 32026
rect 8944 31962 8996 31968
rect 9128 31680 9180 31686
rect 9128 31622 9180 31628
rect 9312 31680 9364 31686
rect 9312 31622 9364 31628
rect 9036 31408 9088 31414
rect 9036 31350 9088 31356
rect 8852 30796 8904 30802
rect 8852 30738 8904 30744
rect 8680 30654 8800 30682
rect 8680 30598 8708 30654
rect 8668 30592 8720 30598
rect 8668 30534 8720 30540
rect 8576 30388 8628 30394
rect 8576 30330 8628 30336
rect 8496 30246 8616 30274
rect 8484 30184 8536 30190
rect 8484 30126 8536 30132
rect 8496 29306 8524 30126
rect 8588 29753 8616 30246
rect 8574 29744 8630 29753
rect 8574 29679 8576 29688
rect 8628 29679 8630 29688
rect 8576 29650 8628 29656
rect 8576 29572 8628 29578
rect 8576 29514 8628 29520
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 8392 29096 8444 29102
rect 8392 29038 8444 29044
rect 8484 27872 8536 27878
rect 8484 27814 8536 27820
rect 8496 26194 8524 27814
rect 8588 27130 8616 29514
rect 8576 27124 8628 27130
rect 8576 27066 8628 27072
rect 8680 27010 8708 30534
rect 8760 29504 8812 29510
rect 8760 29446 8812 29452
rect 8772 29306 8800 29446
rect 8760 29300 8812 29306
rect 8760 29242 8812 29248
rect 8760 28756 8812 28762
rect 8760 28698 8812 28704
rect 8588 26994 8708 27010
rect 8576 26988 8708 26994
rect 8628 26982 8708 26988
rect 8576 26930 8628 26936
rect 8588 26314 8616 26930
rect 8772 26314 8800 28698
rect 8864 27130 8892 30738
rect 8944 30116 8996 30122
rect 8944 30058 8996 30064
rect 8956 29102 8984 30058
rect 8944 29096 8996 29102
rect 8944 29038 8996 29044
rect 9048 28642 9076 31350
rect 9140 29050 9168 31622
rect 9324 30394 9352 31622
rect 9312 30388 9364 30394
rect 9312 30330 9364 30336
rect 9416 30258 9444 32166
rect 9517 32124 9825 32133
rect 9517 32122 9523 32124
rect 9579 32122 9603 32124
rect 9659 32122 9683 32124
rect 9739 32122 9763 32124
rect 9819 32122 9825 32124
rect 9579 32070 9581 32122
rect 9761 32070 9763 32122
rect 9517 32068 9523 32070
rect 9579 32068 9603 32070
rect 9659 32068 9683 32070
rect 9739 32068 9763 32070
rect 9819 32068 9825 32070
rect 9517 32059 9825 32068
rect 9517 31036 9825 31045
rect 9517 31034 9523 31036
rect 9579 31034 9603 31036
rect 9659 31034 9683 31036
rect 9739 31034 9763 31036
rect 9819 31034 9825 31036
rect 9579 30982 9581 31034
rect 9761 30982 9763 31034
rect 9517 30980 9523 30982
rect 9579 30980 9603 30982
rect 9659 30980 9683 30982
rect 9739 30980 9763 30982
rect 9819 30980 9825 30982
rect 9517 30971 9825 30980
rect 9496 30388 9548 30394
rect 9496 30330 9548 30336
rect 9404 30252 9456 30258
rect 9404 30194 9456 30200
rect 9312 30184 9364 30190
rect 9312 30126 9364 30132
rect 9218 29336 9274 29345
rect 9218 29271 9274 29280
rect 9232 29170 9260 29271
rect 9220 29164 9272 29170
rect 9220 29106 9272 29112
rect 9140 29022 9260 29050
rect 9048 28614 9168 28642
rect 9036 28552 9088 28558
rect 9036 28494 9088 28500
rect 9048 28014 9076 28494
rect 9036 28008 9088 28014
rect 9036 27950 9088 27956
rect 8944 27532 8996 27538
rect 8944 27474 8996 27480
rect 8852 27124 8904 27130
rect 8852 27066 8904 27072
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 8760 26308 8812 26314
rect 8760 26250 8812 26256
rect 8496 26166 8616 26194
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 8404 22681 8432 24618
rect 8390 22672 8446 22681
rect 8390 22607 8392 22616
rect 8444 22607 8446 22616
rect 8392 22578 8444 22584
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8404 21554 8432 21830
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8260 21304 8432 21332
rect 8208 21286 8260 21292
rect 8024 21072 8076 21078
rect 8024 21014 8076 21020
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 8208 20868 8260 20874
rect 8208 20810 8260 20816
rect 7576 20760 7678 20788
rect 7742 20760 7880 20788
rect 7576 19378 7604 20760
rect 7742 20618 7770 20760
rect 7803 20700 8111 20709
rect 7803 20698 7809 20700
rect 7865 20698 7889 20700
rect 7945 20698 7969 20700
rect 8025 20698 8049 20700
rect 8105 20698 8111 20700
rect 7865 20646 7867 20698
rect 8047 20646 8049 20698
rect 7803 20644 7809 20646
rect 7865 20644 7889 20646
rect 7945 20644 7969 20646
rect 8025 20644 8049 20646
rect 8105 20644 8111 20646
rect 7803 20635 8111 20644
rect 7668 20590 7770 20618
rect 7932 20596 7984 20602
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7668 19258 7696 20590
rect 7932 20538 7984 20544
rect 7944 20398 7972 20538
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7944 20058 7972 20334
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8220 19938 8248 20810
rect 8404 20466 8432 21304
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8220 19910 8340 19938
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7803 19612 8111 19621
rect 7803 19610 7809 19612
rect 7865 19610 7889 19612
rect 7945 19610 7969 19612
rect 8025 19610 8049 19612
rect 8105 19610 8111 19612
rect 7865 19558 7867 19610
rect 8047 19558 8049 19610
rect 7803 19556 7809 19558
rect 7865 19556 7889 19558
rect 7945 19556 7969 19558
rect 8025 19556 8049 19558
rect 8105 19556 8111 19558
rect 7803 19547 8111 19556
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7576 19230 7696 19258
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7484 12434 7512 18090
rect 7576 17882 7604 19230
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7668 18902 7696 19110
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7668 18737 7696 18838
rect 7654 18728 7710 18737
rect 7654 18663 7710 18672
rect 7760 18612 7788 19450
rect 8220 19378 8248 19790
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8312 19258 8340 19910
rect 8220 19230 8340 19258
rect 7838 19000 7894 19009
rect 7838 18935 7894 18944
rect 7852 18902 7880 18935
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7668 18584 7788 18612
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7562 16552 7618 16561
rect 7562 16487 7618 16496
rect 7576 16114 7604 16487
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7576 13530 7604 13738
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7668 12968 7696 18584
rect 7803 18524 8111 18533
rect 7803 18522 7809 18524
rect 7865 18522 7889 18524
rect 7945 18522 7969 18524
rect 8025 18522 8049 18524
rect 8105 18522 8111 18524
rect 7865 18470 7867 18522
rect 8047 18470 8049 18522
rect 7803 18468 7809 18470
rect 7865 18468 7889 18470
rect 7945 18468 7969 18470
rect 8025 18468 8049 18470
rect 8105 18468 8111 18470
rect 7803 18459 8111 18468
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 8220 17202 8248 19230
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8312 16794 8340 17070
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8404 16674 8432 17818
rect 8312 16646 8432 16674
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 8220 15314 8248 16118
rect 8312 15434 8340 16646
rect 8496 16538 8524 25230
rect 8588 20942 8616 26166
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 8666 24304 8722 24313
rect 8666 24239 8668 24248
rect 8720 24239 8722 24248
rect 8668 24210 8720 24216
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8588 20262 8616 20878
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 18086 8616 18702
rect 8680 18358 8708 24074
rect 8772 22094 8800 24754
rect 8864 23730 8892 27066
rect 8956 26926 8984 27474
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 9048 26858 9076 27950
rect 9036 26852 9088 26858
rect 9036 26794 9088 26800
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8852 23112 8904 23118
rect 8850 23080 8852 23089
rect 8904 23080 8906 23089
rect 8850 23015 8906 23024
rect 8772 22066 8892 22094
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8772 18970 8800 21422
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 17746 8616 18022
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8404 16510 8524 16538
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8404 15348 8432 16510
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8496 15416 8524 16390
rect 8588 15570 8616 17682
rect 8680 17048 8708 18294
rect 8680 17020 8800 17048
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8496 15388 8616 15416
rect 8404 15320 8524 15348
rect 8220 15286 8340 15314
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 8206 15192 8262 15201
rect 8312 15162 8340 15286
rect 8206 15127 8208 15136
rect 8260 15127 8262 15136
rect 8300 15156 8352 15162
rect 8208 15098 8260 15104
rect 8300 15098 8352 15104
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 7840 14068 7892 14074
rect 8220 14056 8248 14214
rect 7840 14010 7892 14016
rect 8128 14028 8248 14056
rect 7852 13870 7880 14010
rect 8128 13938 8156 14028
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8312 13870 8340 14282
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 7668 12940 7788 12968
rect 7484 12406 7696 12434
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 10146 7328 11494
rect 7392 10266 7420 11698
rect 7472 11688 7524 11694
rect 7470 11656 7472 11665
rect 7524 11656 7526 11665
rect 7470 11591 7526 11600
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11354 7512 11494
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7576 11234 7604 12038
rect 7668 11778 7696 12406
rect 7760 12209 7788 12940
rect 8114 12880 8170 12889
rect 8114 12815 8170 12824
rect 8128 12594 8156 12815
rect 8220 12594 8248 13194
rect 8128 12566 8248 12594
rect 7746 12200 7802 12209
rect 7746 12135 7802 12144
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 8220 11914 8248 12566
rect 8220 11886 8340 11914
rect 7668 11750 8248 11778
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7576 11206 8156 11234
rect 7484 10470 7512 11154
rect 7576 10810 7604 11206
rect 8128 11150 8156 11206
rect 7840 11144 7892 11150
rect 7668 11104 7840 11132
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7300 10118 7604 10146
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7194 8528 7250 8537
rect 7194 8463 7250 8472
rect 7208 8430 7236 8463
rect 7392 8430 7420 9590
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7484 9042 7512 9386
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8634 7512 8774
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 3056 1964 3108 1970
rect 3056 1906 3108 1912
rect 5724 1964 5776 1970
rect 5724 1906 5776 1912
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 7196 1964 7248 1970
rect 7196 1906 7248 1912
rect 2663 1660 2971 1669
rect 2663 1658 2669 1660
rect 2725 1658 2749 1660
rect 2805 1658 2829 1660
rect 2885 1658 2909 1660
rect 2965 1658 2971 1660
rect 2725 1606 2727 1658
rect 2907 1606 2909 1658
rect 2663 1604 2669 1606
rect 2725 1604 2749 1606
rect 2805 1604 2829 1606
rect 2885 1604 2909 1606
rect 2965 1604 2971 1606
rect 2663 1595 2971 1604
rect 2136 1352 2188 1358
rect 2056 1312 2136 1340
rect 1584 1284 1636 1290
rect 1584 1226 1636 1232
rect 2056 160 2084 1312
rect 2136 1294 2188 1300
rect 570 0 626 160
rect 1306 0 1362 160
rect 2042 0 2098 160
rect 2778 82 2834 160
rect 3068 82 3096 1906
rect 5736 1562 5764 1906
rect 6090 1660 6398 1669
rect 6090 1658 6096 1660
rect 6152 1658 6176 1660
rect 6232 1658 6256 1660
rect 6312 1658 6336 1660
rect 6392 1658 6398 1660
rect 6152 1606 6154 1658
rect 6334 1606 6336 1658
rect 6090 1604 6096 1606
rect 6152 1604 6176 1606
rect 6232 1604 6256 1606
rect 6312 1604 6336 1606
rect 6392 1604 6398 1606
rect 6090 1595 6398 1604
rect 6472 1562 6500 1906
rect 7208 1562 7236 1906
rect 7392 1834 7420 5170
rect 7576 2774 7604 10118
rect 7668 9654 7696 11104
rect 7840 11086 7892 11092
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7760 10674 7788 10746
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 9042 7880 9318
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8036 9042 8064 9114
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7668 8362 7696 8978
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7668 8090 7696 8298
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 8090 7972 8230
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7668 6254 7696 7278
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 5710 7696 6190
rect 8220 5778 8248 11750
rect 8312 10146 8340 11886
rect 8404 11558 8432 14826
rect 8496 14346 8524 15320
rect 8588 14958 8616 15388
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13530 8524 13806
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8588 13326 8616 14894
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8496 10577 8524 10610
rect 8482 10568 8538 10577
rect 8482 10503 8538 10512
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10266 8432 10406
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8312 10118 8432 10146
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8312 8498 8340 9454
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8404 7818 8432 10118
rect 8588 9110 8616 12922
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8294 8524 8978
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8298 5808 8354 5817
rect 8208 5772 8260 5778
rect 8298 5743 8354 5752
rect 8208 5714 8260 5720
rect 8312 5710 8340 5743
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 7668 5234 7696 5646
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 8404 5234 8432 6938
rect 8496 5914 8524 8230
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8680 4554 8708 16526
rect 8772 15366 8800 17020
rect 8864 16590 8892 22066
rect 8956 21486 8984 24550
rect 9048 22250 9076 26794
rect 9140 24206 9168 28614
rect 9232 28529 9260 29022
rect 9324 28694 9352 30126
rect 9508 30036 9536 30330
rect 9416 30008 9536 30036
rect 9312 28688 9364 28694
rect 9312 28630 9364 28636
rect 9218 28520 9274 28529
rect 9416 28506 9444 30008
rect 9517 29948 9825 29957
rect 9517 29946 9523 29948
rect 9579 29946 9603 29948
rect 9659 29946 9683 29948
rect 9739 29946 9763 29948
rect 9819 29946 9825 29948
rect 9579 29894 9581 29946
rect 9761 29894 9763 29946
rect 9517 29892 9523 29894
rect 9579 29892 9603 29894
rect 9659 29892 9683 29894
rect 9739 29892 9763 29894
rect 9819 29892 9825 29894
rect 9517 29883 9825 29892
rect 9586 29744 9642 29753
rect 9586 29679 9642 29688
rect 9600 29050 9628 29679
rect 9876 29306 9904 32506
rect 10152 31346 10180 33254
rect 10336 32434 10364 33798
rect 10324 32428 10376 32434
rect 10324 32370 10376 32376
rect 10428 32026 10456 34598
rect 10888 34610 10916 36094
rect 10966 36071 11022 36080
rect 11072 35154 11100 36722
rect 12176 36378 12204 36722
rect 12268 36650 12296 37674
rect 12360 37126 12388 38830
rect 12728 38554 12756 38898
rect 12808 38752 12860 38758
rect 12808 38694 12860 38700
rect 12716 38548 12768 38554
rect 12716 38490 12768 38496
rect 12716 38412 12768 38418
rect 12716 38354 12768 38360
rect 12624 38344 12676 38350
rect 12624 38286 12676 38292
rect 12636 38010 12664 38286
rect 12624 38004 12676 38010
rect 12624 37946 12676 37952
rect 12624 37800 12676 37806
rect 12624 37742 12676 37748
rect 12636 37466 12664 37742
rect 12624 37460 12676 37466
rect 12624 37402 12676 37408
rect 12532 37256 12584 37262
rect 12532 37198 12584 37204
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 12256 36644 12308 36650
rect 12256 36586 12308 36592
rect 12348 36644 12400 36650
rect 12348 36586 12400 36592
rect 12360 36378 12388 36586
rect 12440 36576 12492 36582
rect 12440 36518 12492 36524
rect 12164 36372 12216 36378
rect 12164 36314 12216 36320
rect 12348 36372 12400 36378
rect 12348 36314 12400 36320
rect 11796 36168 11848 36174
rect 11796 36110 11848 36116
rect 12164 36168 12216 36174
rect 12164 36110 12216 36116
rect 11230 35932 11538 35941
rect 11230 35930 11236 35932
rect 11292 35930 11316 35932
rect 11372 35930 11396 35932
rect 11452 35930 11476 35932
rect 11532 35930 11538 35932
rect 11292 35878 11294 35930
rect 11474 35878 11476 35930
rect 11230 35876 11236 35878
rect 11292 35876 11316 35878
rect 11372 35876 11396 35878
rect 11452 35876 11476 35878
rect 11532 35876 11538 35878
rect 11230 35867 11538 35876
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 11520 35148 11572 35154
rect 11572 35108 11652 35136
rect 11520 35090 11572 35096
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 10980 34746 11008 35022
rect 11152 35012 11204 35018
rect 11152 34954 11204 34960
rect 10968 34740 11020 34746
rect 10968 34682 11020 34688
rect 10690 34575 10746 34584
rect 10876 34604 10928 34610
rect 10600 34546 10652 34552
rect 10508 34536 10560 34542
rect 10508 34478 10560 34484
rect 10520 34202 10548 34478
rect 10508 34196 10560 34202
rect 10508 34138 10560 34144
rect 10508 33856 10560 33862
rect 10508 33798 10560 33804
rect 10416 32020 10468 32026
rect 10416 31962 10468 31968
rect 10520 31906 10548 33798
rect 10244 31878 10548 31906
rect 10140 31340 10192 31346
rect 10140 31282 10192 31288
rect 10152 30598 10180 31282
rect 10140 30592 10192 30598
rect 10140 30534 10192 30540
rect 10140 30184 10192 30190
rect 10140 30126 10192 30132
rect 9956 30048 10008 30054
rect 9956 29990 10008 29996
rect 9968 29782 9996 29990
rect 10048 29844 10100 29850
rect 10048 29786 10100 29792
rect 9956 29776 10008 29782
rect 9956 29718 10008 29724
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9864 29300 9916 29306
rect 9864 29242 9916 29248
rect 9864 29096 9916 29102
rect 9784 29056 9864 29084
rect 9784 29050 9812 29056
rect 9600 29022 9812 29050
rect 9864 29038 9916 29044
rect 9517 28860 9825 28869
rect 9517 28858 9523 28860
rect 9579 28858 9603 28860
rect 9659 28858 9683 28860
rect 9739 28858 9763 28860
rect 9819 28858 9825 28860
rect 9579 28806 9581 28858
rect 9761 28806 9763 28858
rect 9517 28804 9523 28806
rect 9579 28804 9603 28806
rect 9659 28804 9683 28806
rect 9739 28804 9763 28806
rect 9819 28804 9825 28806
rect 9517 28795 9825 28804
rect 9588 28756 9640 28762
rect 9588 28698 9640 28704
rect 9600 28642 9628 28698
rect 9968 28694 9996 29446
rect 9956 28688 10008 28694
rect 9496 28620 9548 28626
rect 9600 28614 9720 28642
rect 9956 28630 10008 28636
rect 9496 28562 9548 28568
rect 9218 28455 9274 28464
rect 9324 28478 9444 28506
rect 9232 27470 9260 28455
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 9232 24750 9260 25774
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9232 23526 9260 24686
rect 9324 24206 9352 28478
rect 9508 28370 9536 28562
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9416 28342 9536 28370
rect 9416 28014 9444 28342
rect 9600 28218 9628 28494
rect 9588 28212 9640 28218
rect 9588 28154 9640 28160
rect 9600 28121 9628 28154
rect 9586 28112 9642 28121
rect 9586 28047 9642 28056
rect 9404 28008 9456 28014
rect 9692 27962 9720 28614
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 9968 28098 9996 28154
rect 9784 28082 9996 28098
rect 9772 28076 9996 28082
rect 9824 28070 9996 28076
rect 9772 28018 9824 28024
rect 9404 27950 9456 27956
rect 9600 27934 9720 27962
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 9600 27860 9628 27934
rect 9416 27832 9628 27860
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9416 24018 9444 27832
rect 9517 27772 9825 27781
rect 9517 27770 9523 27772
rect 9579 27770 9603 27772
rect 9659 27770 9683 27772
rect 9739 27770 9763 27772
rect 9819 27770 9825 27772
rect 9579 27718 9581 27770
rect 9761 27718 9763 27770
rect 9517 27716 9523 27718
rect 9579 27716 9603 27718
rect 9659 27716 9683 27718
rect 9739 27716 9763 27718
rect 9819 27716 9825 27718
rect 9517 27707 9825 27716
rect 9876 27674 9904 27950
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9862 27432 9918 27441
rect 9862 27367 9918 27376
rect 9876 26926 9904 27367
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9517 26684 9825 26693
rect 9517 26682 9523 26684
rect 9579 26682 9603 26684
rect 9659 26682 9683 26684
rect 9739 26682 9763 26684
rect 9819 26682 9825 26684
rect 9579 26630 9581 26682
rect 9761 26630 9763 26682
rect 9517 26628 9523 26630
rect 9579 26628 9603 26630
rect 9659 26628 9683 26630
rect 9739 26628 9763 26630
rect 9819 26628 9825 26630
rect 9517 26619 9825 26628
rect 9876 26450 9904 26862
rect 9864 26444 9916 26450
rect 9864 26386 9916 26392
rect 9517 25596 9825 25605
rect 9517 25594 9523 25596
rect 9579 25594 9603 25596
rect 9659 25594 9683 25596
rect 9739 25594 9763 25596
rect 9819 25594 9825 25596
rect 9579 25542 9581 25594
rect 9761 25542 9763 25594
rect 9517 25540 9523 25542
rect 9579 25540 9603 25542
rect 9659 25540 9683 25542
rect 9739 25540 9763 25542
rect 9819 25540 9825 25542
rect 9517 25531 9825 25540
rect 9496 25356 9548 25362
rect 9496 25298 9548 25304
rect 9508 24954 9536 25298
rect 9968 25294 9996 28070
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9876 24954 9904 25230
rect 9496 24948 9548 24954
rect 9496 24890 9548 24896
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9876 24614 9904 24890
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9517 24508 9825 24517
rect 9517 24506 9523 24508
rect 9579 24506 9603 24508
rect 9659 24506 9683 24508
rect 9739 24506 9763 24508
rect 9819 24506 9825 24508
rect 9579 24454 9581 24506
rect 9761 24454 9763 24506
rect 9517 24452 9523 24454
rect 9579 24452 9603 24454
rect 9659 24452 9683 24454
rect 9739 24452 9763 24454
rect 9819 24452 9825 24454
rect 9517 24443 9825 24452
rect 9494 24304 9550 24313
rect 9494 24239 9550 24248
rect 9324 23990 9444 24018
rect 9220 23520 9272 23526
rect 9220 23462 9272 23468
rect 9128 22432 9180 22438
rect 9180 22392 9260 22420
rect 9128 22374 9180 22380
rect 9048 22222 9168 22250
rect 9036 22160 9088 22166
rect 9036 22102 9088 22108
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8942 20904 8998 20913
rect 8942 20839 8998 20848
rect 8956 19922 8984 20839
rect 9048 19938 9076 22102
rect 9140 21486 9168 22222
rect 9232 21554 9260 22392
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 9324 20262 9352 23990
rect 9508 23576 9536 24239
rect 9416 23548 9536 23576
rect 9416 23186 9444 23548
rect 9517 23420 9825 23429
rect 9517 23418 9523 23420
rect 9579 23418 9603 23420
rect 9659 23418 9683 23420
rect 9739 23418 9763 23420
rect 9819 23418 9825 23420
rect 9579 23366 9581 23418
rect 9761 23366 9763 23418
rect 9517 23364 9523 23366
rect 9579 23364 9603 23366
rect 9659 23364 9683 23366
rect 9739 23364 9763 23366
rect 9819 23364 9825 23366
rect 9517 23355 9825 23364
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9416 22642 9444 23122
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 20534 9444 22374
rect 9517 22332 9825 22341
rect 9517 22330 9523 22332
rect 9579 22330 9603 22332
rect 9659 22330 9683 22332
rect 9739 22330 9763 22332
rect 9819 22330 9825 22332
rect 9579 22278 9581 22330
rect 9761 22278 9763 22330
rect 9517 22276 9523 22278
rect 9579 22276 9603 22278
rect 9659 22276 9683 22278
rect 9739 22276 9763 22278
rect 9819 22276 9825 22278
rect 9517 22267 9825 22276
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9784 21729 9812 22034
rect 9862 21992 9918 22001
rect 9862 21927 9918 21936
rect 9770 21720 9826 21729
rect 9876 21690 9904 21927
rect 9968 21876 9996 25230
rect 10060 21978 10088 29786
rect 10152 29646 10180 30126
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10152 27538 10180 29582
rect 10140 27532 10192 27538
rect 10140 27474 10192 27480
rect 10140 27396 10192 27402
rect 10140 27338 10192 27344
rect 10152 26353 10180 27338
rect 10244 26382 10272 31878
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10324 30864 10376 30870
rect 10324 30806 10376 30812
rect 10336 28762 10364 30806
rect 10324 28756 10376 28762
rect 10324 28698 10376 28704
rect 10428 28626 10456 31078
rect 10508 30728 10560 30734
rect 10508 30670 10560 30676
rect 10416 28620 10468 28626
rect 10416 28562 10468 28568
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10336 28218 10364 28494
rect 10520 28218 10548 30670
rect 10324 28212 10376 28218
rect 10324 28154 10376 28160
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10324 27532 10376 27538
rect 10324 27474 10376 27480
rect 10232 26376 10284 26382
rect 10138 26344 10194 26353
rect 10232 26318 10284 26324
rect 10138 26279 10194 26288
rect 10244 25906 10272 26318
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10232 23792 10284 23798
rect 10232 23734 10284 23740
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10152 22098 10180 23462
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10060 21950 10180 21978
rect 9968 21848 10088 21876
rect 9770 21655 9826 21664
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9517 21244 9825 21253
rect 9517 21242 9523 21244
rect 9579 21242 9603 21244
rect 9659 21242 9683 21244
rect 9739 21242 9763 21244
rect 9819 21242 9825 21244
rect 9579 21190 9581 21242
rect 9761 21190 9763 21242
rect 9517 21188 9523 21190
rect 9579 21188 9603 21190
rect 9659 21188 9683 21190
rect 9739 21188 9763 21190
rect 9819 21188 9825 21190
rect 9517 21179 9825 21188
rect 9772 20936 9824 20942
rect 9824 20896 9904 20924
rect 9772 20878 9824 20884
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9692 20534 9720 20810
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9232 20058 9260 20198
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 8944 19916 8996 19922
rect 9048 19910 9260 19938
rect 8944 19858 8996 19864
rect 8956 19258 8984 19858
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9034 19544 9090 19553
rect 9034 19479 9036 19488
rect 9088 19479 9090 19488
rect 9036 19450 9088 19456
rect 8956 19230 9076 19258
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8956 16726 8984 19110
rect 8944 16720 8996 16726
rect 8944 16662 8996 16668
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8942 16144 8998 16153
rect 8942 16079 8944 16088
rect 8996 16079 8998 16088
rect 8944 16050 8996 16056
rect 9048 15960 9076 19230
rect 8864 15932 9076 15960
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8864 14414 8892 15932
rect 9140 15910 9168 19790
rect 9232 17882 9260 19910
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9324 17338 9352 19654
rect 9416 19242 9444 20334
rect 9517 20156 9825 20165
rect 9517 20154 9523 20156
rect 9579 20154 9603 20156
rect 9659 20154 9683 20156
rect 9739 20154 9763 20156
rect 9819 20154 9825 20156
rect 9579 20102 9581 20154
rect 9761 20102 9763 20154
rect 9517 20100 9523 20102
rect 9579 20100 9603 20102
rect 9659 20100 9683 20102
rect 9739 20100 9763 20102
rect 9819 20100 9825 20102
rect 9517 20091 9825 20100
rect 9876 20040 9904 20896
rect 9692 20012 9904 20040
rect 9954 20088 10010 20097
rect 10060 20074 10088 21848
rect 10152 20097 10180 21950
rect 10010 20046 10088 20074
rect 10138 20088 10194 20097
rect 9954 20023 10010 20032
rect 10138 20023 10194 20032
rect 9692 19334 9720 20012
rect 10244 19938 10272 23734
rect 10336 22778 10364 27474
rect 10612 25498 10640 34546
rect 10704 33114 10732 34575
rect 10876 34546 10928 34552
rect 11060 34604 11112 34610
rect 11060 34546 11112 34552
rect 11072 34490 11100 34546
rect 10888 34462 11100 34490
rect 10784 33584 10836 33590
rect 10784 33526 10836 33532
rect 10692 33108 10744 33114
rect 10692 33050 10744 33056
rect 10796 32026 10824 33526
rect 10888 32978 10916 34462
rect 11164 34354 11192 34954
rect 11230 34844 11538 34853
rect 11230 34842 11236 34844
rect 11292 34842 11316 34844
rect 11372 34842 11396 34844
rect 11452 34842 11476 34844
rect 11532 34842 11538 34844
rect 11292 34790 11294 34842
rect 11474 34790 11476 34842
rect 11230 34788 11236 34790
rect 11292 34788 11316 34790
rect 11372 34788 11396 34790
rect 11452 34788 11476 34790
rect 11532 34788 11538 34790
rect 11230 34779 11538 34788
rect 11072 34326 11192 34354
rect 10876 32972 10928 32978
rect 10876 32914 10928 32920
rect 11072 32858 11100 34326
rect 11624 34066 11652 35108
rect 11612 34060 11664 34066
rect 11612 34002 11664 34008
rect 11520 33992 11572 33998
rect 11518 33960 11520 33969
rect 11572 33960 11574 33969
rect 11624 33930 11652 34002
rect 11808 33998 11836 36110
rect 12072 36032 12124 36038
rect 11900 35992 12072 36020
rect 11900 35698 11928 35992
rect 12072 35974 12124 35980
rect 11888 35692 11940 35698
rect 12072 35692 12124 35698
rect 11888 35634 11940 35640
rect 11992 35652 12072 35680
rect 11992 34762 12020 35652
rect 12072 35634 12124 35640
rect 12176 35086 12204 36110
rect 12452 35766 12480 36518
rect 12440 35760 12492 35766
rect 12440 35702 12492 35708
rect 12544 35193 12572 37198
rect 12624 36916 12676 36922
rect 12728 36904 12756 38354
rect 12820 38214 12848 38694
rect 12944 38652 13252 38661
rect 12944 38650 12950 38652
rect 13006 38650 13030 38652
rect 13086 38650 13110 38652
rect 13166 38650 13190 38652
rect 13246 38650 13252 38652
rect 13006 38598 13008 38650
rect 13188 38598 13190 38650
rect 12944 38596 12950 38598
rect 13006 38596 13030 38598
rect 13086 38596 13110 38598
rect 13166 38596 13190 38598
rect 13246 38596 13252 38598
rect 12944 38587 13252 38596
rect 13280 38554 13308 39374
rect 13544 39364 13596 39370
rect 13544 39306 13596 39312
rect 13912 39364 13964 39370
rect 13912 39306 13964 39312
rect 13556 39098 13584 39306
rect 13544 39092 13596 39098
rect 13544 39034 13596 39040
rect 13924 39001 13952 39306
rect 13910 38992 13966 39001
rect 13360 38956 13412 38962
rect 13910 38927 13966 38936
rect 14004 38956 14056 38962
rect 13360 38898 13412 38904
rect 14004 38898 14056 38904
rect 13268 38548 13320 38554
rect 13268 38490 13320 38496
rect 12808 38208 12860 38214
rect 12808 38150 12860 38156
rect 13268 38208 13320 38214
rect 13268 38150 13320 38156
rect 12676 36876 12756 36904
rect 12624 36858 12676 36864
rect 12716 36780 12768 36786
rect 12716 36722 12768 36728
rect 12728 36378 12756 36722
rect 12716 36372 12768 36378
rect 12716 36314 12768 36320
rect 12820 36258 12848 38150
rect 13280 37942 13308 38150
rect 13268 37936 13320 37942
rect 13268 37878 13320 37884
rect 13372 37670 13400 38898
rect 13544 38888 13596 38894
rect 13544 38830 13596 38836
rect 13452 38344 13504 38350
rect 13452 38286 13504 38292
rect 13556 38298 13584 38830
rect 13820 38820 13872 38826
rect 13820 38762 13872 38768
rect 13636 38752 13688 38758
rect 13636 38694 13688 38700
rect 13648 38457 13676 38694
rect 13634 38448 13690 38457
rect 13634 38383 13690 38392
rect 13832 38350 13860 38762
rect 13820 38344 13872 38350
rect 13360 37664 13412 37670
rect 13360 37606 13412 37612
rect 12944 37564 13252 37573
rect 12944 37562 12950 37564
rect 13006 37562 13030 37564
rect 13086 37562 13110 37564
rect 13166 37562 13190 37564
rect 13246 37562 13252 37564
rect 13006 37510 13008 37562
rect 13188 37510 13190 37562
rect 12944 37508 12950 37510
rect 13006 37508 13030 37510
rect 13086 37508 13110 37510
rect 13166 37508 13190 37510
rect 13246 37508 13252 37510
rect 12944 37499 13252 37508
rect 13084 37256 13136 37262
rect 13082 37224 13084 37233
rect 13360 37256 13412 37262
rect 13136 37224 13138 37233
rect 13360 37198 13412 37204
rect 13082 37159 13138 37168
rect 13084 37120 13136 37126
rect 13084 37062 13136 37068
rect 13096 36922 13124 37062
rect 13084 36916 13136 36922
rect 13084 36858 13136 36864
rect 13268 36712 13320 36718
rect 13268 36654 13320 36660
rect 12944 36476 13252 36485
rect 12944 36474 12950 36476
rect 13006 36474 13030 36476
rect 13086 36474 13110 36476
rect 13166 36474 13190 36476
rect 13246 36474 13252 36476
rect 13006 36422 13008 36474
rect 13188 36422 13190 36474
rect 12944 36420 12950 36422
rect 13006 36420 13030 36422
rect 13086 36420 13110 36422
rect 13166 36420 13190 36422
rect 13246 36420 13252 36422
rect 12944 36411 13252 36420
rect 13280 36281 13308 36654
rect 13372 36378 13400 37198
rect 13464 36689 13492 38286
rect 13556 38270 13676 38298
rect 13820 38286 13872 38292
rect 13544 37868 13596 37874
rect 13544 37810 13596 37816
rect 13556 37466 13584 37810
rect 13544 37460 13596 37466
rect 13544 37402 13596 37408
rect 13648 36938 13676 38270
rect 13820 38208 13872 38214
rect 13820 38150 13872 38156
rect 13832 37913 13860 38150
rect 14016 37942 14044 38898
rect 14188 38752 14240 38758
rect 14188 38694 14240 38700
rect 14200 38593 14228 38694
rect 14186 38584 14242 38593
rect 14186 38519 14242 38528
rect 14004 37936 14056 37942
rect 13818 37904 13874 37913
rect 14004 37878 14056 37884
rect 13818 37839 13874 37848
rect 14004 37800 14056 37806
rect 14004 37742 14056 37748
rect 13728 37664 13780 37670
rect 13728 37606 13780 37612
rect 13556 36910 13676 36938
rect 13450 36680 13506 36689
rect 13450 36615 13506 36624
rect 13556 36530 13584 36910
rect 13636 36848 13688 36854
rect 13740 36825 13768 37606
rect 14016 37369 14044 37742
rect 14002 37360 14058 37369
rect 14002 37295 14058 37304
rect 13636 36790 13688 36796
rect 13726 36816 13782 36825
rect 13464 36502 13584 36530
rect 13360 36372 13412 36378
rect 13360 36314 13412 36320
rect 12636 36230 12848 36258
rect 13266 36272 13322 36281
rect 12530 35184 12586 35193
rect 12530 35119 12586 35128
rect 12164 35080 12216 35086
rect 12164 35022 12216 35028
rect 12348 34944 12400 34950
rect 11900 34734 12020 34762
rect 12084 34904 12348 34932
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 11518 33895 11574 33904
rect 11612 33924 11664 33930
rect 11612 33866 11664 33872
rect 11230 33756 11538 33765
rect 11230 33754 11236 33756
rect 11292 33754 11316 33756
rect 11372 33754 11396 33756
rect 11452 33754 11476 33756
rect 11532 33754 11538 33756
rect 11292 33702 11294 33754
rect 11474 33702 11476 33754
rect 11230 33700 11236 33702
rect 11292 33700 11316 33702
rect 11372 33700 11396 33702
rect 11452 33700 11476 33702
rect 11532 33700 11538 33702
rect 11230 33691 11538 33700
rect 11624 33454 11652 33866
rect 11796 33516 11848 33522
rect 11796 33458 11848 33464
rect 11612 33448 11664 33454
rect 11612 33390 11664 33396
rect 10888 32830 11100 32858
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 10888 32314 10916 32830
rect 11060 32768 11112 32774
rect 11060 32710 11112 32716
rect 11072 32434 11100 32710
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 10888 32286 11008 32314
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10784 31816 10836 31822
rect 10784 31758 10836 31764
rect 10980 31770 11008 32286
rect 11072 31929 11100 32370
rect 11058 31920 11114 31929
rect 11058 31855 11114 31864
rect 10796 31482 10824 31758
rect 10876 31748 10928 31754
rect 10980 31742 11100 31770
rect 10876 31690 10928 31696
rect 10888 31482 10916 31690
rect 10784 31476 10836 31482
rect 10784 31418 10836 31424
rect 10876 31476 10928 31482
rect 10876 31418 10928 31424
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 10796 30025 10824 31078
rect 10888 30938 10916 31282
rect 10876 30932 10928 30938
rect 10876 30874 10928 30880
rect 11072 30784 11100 31742
rect 10888 30756 11100 30784
rect 10888 30394 10916 30756
rect 11060 30660 11112 30666
rect 11060 30602 11112 30608
rect 10876 30388 10928 30394
rect 10876 30330 10928 30336
rect 10876 30252 10928 30258
rect 10876 30194 10928 30200
rect 10782 30016 10838 30025
rect 10782 29951 10838 29960
rect 10690 29880 10746 29889
rect 10690 29815 10692 29824
rect 10744 29815 10746 29824
rect 10784 29844 10836 29850
rect 10692 29786 10744 29792
rect 10784 29786 10836 29792
rect 10692 28416 10744 28422
rect 10692 28358 10744 28364
rect 10704 27062 10732 28358
rect 10692 27056 10744 27062
rect 10692 26998 10744 27004
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10414 25120 10470 25129
rect 10414 25055 10470 25064
rect 10428 24818 10456 25055
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10336 22166 10364 22714
rect 10324 22160 10376 22166
rect 10324 22102 10376 22108
rect 10520 22098 10548 22918
rect 10508 22092 10560 22098
rect 10428 22052 10508 22080
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 9874 19922 10272 19938
rect 9862 19916 10272 19922
rect 9914 19910 10272 19916
rect 9862 19858 9914 19864
rect 9956 19848 10008 19854
rect 10008 19796 10021 19836
rect 9956 19790 10021 19796
rect 9968 19774 10021 19790
rect 9862 19680 9918 19689
rect 9968 19666 9996 19774
rect 10138 19680 10194 19689
rect 9968 19638 10138 19666
rect 9862 19615 9918 19624
rect 10138 19615 10194 19624
rect 9876 19530 9904 19615
rect 10046 19544 10102 19553
rect 9876 19502 9996 19530
rect 9692 19306 9904 19334
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9416 18222 9444 19178
rect 9517 19068 9825 19077
rect 9517 19066 9523 19068
rect 9579 19066 9603 19068
rect 9659 19066 9683 19068
rect 9739 19066 9763 19068
rect 9819 19066 9825 19068
rect 9579 19014 9581 19066
rect 9761 19014 9763 19066
rect 9517 19012 9523 19014
rect 9579 19012 9603 19014
rect 9659 19012 9683 19014
rect 9739 19012 9763 19014
rect 9819 19012 9825 19014
rect 9517 19003 9825 19012
rect 9680 18896 9732 18902
rect 9586 18864 9642 18873
rect 9680 18838 9732 18844
rect 9586 18799 9642 18808
rect 9600 18290 9628 18799
rect 9692 18737 9720 18838
rect 9876 18766 9904 19306
rect 9968 19242 9996 19502
rect 10046 19479 10102 19488
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9864 18760 9916 18766
rect 9678 18728 9734 18737
rect 9864 18702 9916 18708
rect 9678 18663 9734 18672
rect 10060 18578 10088 19479
rect 9876 18550 10088 18578
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9416 17134 9444 18022
rect 9517 17980 9825 17989
rect 9517 17978 9523 17980
rect 9579 17978 9603 17980
rect 9659 17978 9683 17980
rect 9739 17978 9763 17980
rect 9819 17978 9825 17980
rect 9579 17926 9581 17978
rect 9761 17926 9763 17978
rect 9517 17924 9523 17926
rect 9579 17924 9603 17926
rect 9659 17924 9683 17926
rect 9739 17924 9763 17926
rect 9819 17924 9825 17926
rect 9517 17915 9825 17924
rect 9678 17776 9734 17785
rect 9678 17711 9734 17720
rect 9692 17678 9720 17711
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9404 17128 9456 17134
rect 9692 17105 9720 17614
rect 9876 17202 9904 18550
rect 10152 18442 10180 19615
rect 9968 18414 10180 18442
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9404 17070 9456 17076
rect 9678 17096 9734 17105
rect 9678 17031 9734 17040
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 9218 16552 9274 16561
rect 9218 16487 9274 16496
rect 9588 16516 9640 16522
rect 9128 15904 9180 15910
rect 8956 15864 9128 15892
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 14006 8892 14214
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8772 11354 8800 12310
rect 8864 11830 8892 13262
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8850 11656 8906 11665
rect 8850 11591 8906 11600
rect 8864 11354 8892 11591
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8956 11234 8984 15864
rect 9128 15846 9180 15852
rect 9232 15502 9260 16487
rect 9588 16458 9640 16464
rect 9310 16144 9366 16153
rect 9310 16079 9366 16088
rect 9220 15496 9272 15502
rect 9048 15444 9220 15450
rect 9048 15438 9272 15444
rect 9048 15422 9260 15438
rect 9048 14890 9076 15422
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9036 14000 9088 14006
rect 9034 13968 9036 13977
rect 9088 13968 9090 13977
rect 9034 13903 9090 13912
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 11370 9076 13670
rect 9140 12170 9168 14554
rect 9232 13852 9260 15302
rect 9324 14074 9352 16079
rect 9600 16046 9628 16458
rect 9876 16402 9904 17138
rect 9968 16810 9996 18414
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10152 18057 10180 18158
rect 10138 18048 10194 18057
rect 10138 17983 10194 17992
rect 10048 16992 10100 16998
rect 10100 16952 10180 16980
rect 10048 16934 10100 16940
rect 10152 16833 10180 16952
rect 10138 16824 10194 16833
rect 9968 16782 10088 16810
rect 9954 16416 10010 16425
rect 9876 16374 9954 16402
rect 9954 16351 10010 16360
rect 9588 16040 9640 16046
rect 9416 16000 9588 16028
rect 9416 14618 9444 16000
rect 9588 15982 9640 15988
rect 9772 16040 9824 16046
rect 9824 16000 9996 16028
rect 9772 15982 9824 15988
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 9968 15706 9996 16000
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 10060 15586 10088 16782
rect 10138 16759 10194 16768
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 9968 15558 10088 15586
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9784 14958 9812 15438
rect 9772 14952 9824 14958
rect 9824 14912 9904 14940
rect 9772 14894 9824 14900
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9600 14346 9628 14486
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9784 13938 9812 14350
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9232 13824 9352 13852
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9232 11830 9260 12038
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9048 11342 9168 11370
rect 8956 11206 9076 11234
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10062 8800 10950
rect 8850 10704 8906 10713
rect 8850 10639 8906 10648
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 8090 8800 8910
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 7576 2746 7696 2774
rect 7668 2106 7696 2746
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 8864 2106 8892 10639
rect 8956 9450 8984 11018
rect 8944 9444 8996 9450
rect 8944 9386 8996 9392
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 8852 2100 8904 2106
rect 8852 2042 8904 2048
rect 8956 2038 8984 9046
rect 9048 7410 9076 11206
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 6769 9076 7346
rect 9034 6760 9090 6769
rect 9034 6695 9090 6704
rect 9048 6322 9076 6695
rect 9140 6644 9168 11342
rect 9324 11150 9352 13824
rect 9416 13530 9444 13874
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9416 12850 9444 13194
rect 9876 13190 9904 14912
rect 9968 13977 9996 15558
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14006 10088 14758
rect 10048 14000 10100 14006
rect 9954 13968 10010 13977
rect 10048 13942 10100 13948
rect 9954 13903 10010 13912
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 10060 12850 10088 13330
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 9994 9352 10610
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9416 9058 9444 12786
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 9864 12436 9916 12442
rect 10152 12434 10180 16526
rect 10244 14822 10272 19910
rect 10336 19378 10364 21830
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 17082 10364 18634
rect 10428 17921 10456 22052
rect 10612 22094 10640 25434
rect 10704 24188 10732 25774
rect 10796 25498 10824 29786
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 10784 24200 10836 24206
rect 10704 24160 10784 24188
rect 10784 24142 10836 24148
rect 10796 23798 10824 24142
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10888 23118 10916 30194
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10980 28506 11008 29990
rect 11072 29238 11100 30602
rect 11164 30122 11192 32846
rect 11230 32668 11538 32677
rect 11230 32666 11236 32668
rect 11292 32666 11316 32668
rect 11372 32666 11396 32668
rect 11452 32666 11476 32668
rect 11532 32666 11538 32668
rect 11292 32614 11294 32666
rect 11474 32614 11476 32666
rect 11230 32612 11236 32614
rect 11292 32612 11316 32614
rect 11372 32612 11396 32614
rect 11452 32612 11476 32614
rect 11532 32612 11538 32614
rect 11230 32603 11538 32612
rect 11520 32360 11572 32366
rect 11624 32348 11652 33390
rect 11808 33114 11836 33458
rect 11796 33108 11848 33114
rect 11796 33050 11848 33056
rect 11900 32960 11928 34734
rect 11980 34672 12032 34678
rect 11980 34614 12032 34620
rect 11572 32320 11652 32348
rect 11716 32932 11928 32960
rect 11520 32302 11572 32308
rect 11518 31920 11574 31929
rect 11518 31855 11574 31864
rect 11532 31822 11560 31855
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11612 31816 11664 31822
rect 11612 31758 11664 31764
rect 11230 31580 11538 31589
rect 11230 31578 11236 31580
rect 11292 31578 11316 31580
rect 11372 31578 11396 31580
rect 11452 31578 11476 31580
rect 11532 31578 11538 31580
rect 11292 31526 11294 31578
rect 11474 31526 11476 31578
rect 11230 31524 11236 31526
rect 11292 31524 11316 31526
rect 11372 31524 11396 31526
rect 11452 31524 11476 31526
rect 11532 31524 11538 31526
rect 11230 31515 11538 31524
rect 11244 31272 11296 31278
rect 11244 31214 11296 31220
rect 11256 30841 11284 31214
rect 11242 30832 11298 30841
rect 11242 30767 11298 30776
rect 11230 30492 11538 30501
rect 11230 30490 11236 30492
rect 11292 30490 11316 30492
rect 11372 30490 11396 30492
rect 11452 30490 11476 30492
rect 11532 30490 11538 30492
rect 11292 30438 11294 30490
rect 11474 30438 11476 30490
rect 11230 30436 11236 30438
rect 11292 30436 11316 30438
rect 11372 30436 11396 30438
rect 11452 30436 11476 30438
rect 11532 30436 11538 30438
rect 11230 30427 11538 30436
rect 11336 30320 11388 30326
rect 11624 30297 11652 31758
rect 11336 30262 11388 30268
rect 11610 30288 11666 30297
rect 11152 30116 11204 30122
rect 11152 30058 11204 30064
rect 11244 30048 11296 30054
rect 11150 30016 11206 30025
rect 11348 30025 11376 30262
rect 11520 30252 11572 30258
rect 11610 30223 11666 30232
rect 11520 30194 11572 30200
rect 11532 30138 11560 30194
rect 11532 30110 11652 30138
rect 11244 29990 11296 29996
rect 11334 30016 11390 30025
rect 11150 29951 11206 29960
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 11072 28801 11100 28902
rect 11058 28792 11114 28801
rect 11058 28727 11114 28736
rect 11058 28520 11114 28529
rect 10980 28478 11058 28506
rect 11058 28455 11114 28464
rect 11164 28200 11192 29951
rect 11256 29753 11284 29990
rect 11334 29951 11390 29960
rect 11426 29880 11482 29889
rect 11426 29815 11482 29824
rect 11336 29776 11388 29782
rect 11242 29744 11298 29753
rect 11336 29718 11388 29724
rect 11242 29679 11298 29688
rect 11244 29640 11296 29646
rect 11242 29608 11244 29617
rect 11296 29608 11298 29617
rect 11348 29578 11376 29718
rect 11440 29646 11468 29815
rect 11428 29640 11480 29646
rect 11428 29582 11480 29588
rect 11242 29543 11298 29552
rect 11336 29572 11388 29578
rect 11336 29514 11388 29520
rect 11230 29404 11538 29413
rect 11230 29402 11236 29404
rect 11292 29402 11316 29404
rect 11372 29402 11396 29404
rect 11452 29402 11476 29404
rect 11532 29402 11538 29404
rect 11292 29350 11294 29402
rect 11474 29350 11476 29402
rect 11230 29348 11236 29350
rect 11292 29348 11316 29350
rect 11372 29348 11396 29350
rect 11452 29348 11476 29350
rect 11532 29348 11538 29350
rect 11230 29339 11538 29348
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11256 29186 11284 29242
rect 11624 29186 11652 30110
rect 11256 29158 11652 29186
rect 11256 29034 11284 29158
rect 11610 29064 11666 29073
rect 11244 29028 11296 29034
rect 11244 28970 11296 28976
rect 11520 29028 11572 29034
rect 11610 28999 11666 29008
rect 11520 28970 11572 28976
rect 11532 28422 11560 28970
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11230 28316 11538 28325
rect 11230 28314 11236 28316
rect 11292 28314 11316 28316
rect 11372 28314 11396 28316
rect 11452 28314 11476 28316
rect 11532 28314 11538 28316
rect 11292 28262 11294 28314
rect 11474 28262 11476 28314
rect 11230 28260 11236 28262
rect 11292 28260 11316 28262
rect 11372 28260 11396 28262
rect 11452 28260 11476 28262
rect 11532 28260 11538 28262
rect 11230 28251 11538 28260
rect 10980 28172 11192 28200
rect 10980 27062 11008 28172
rect 11520 28008 11572 28014
rect 11520 27950 11572 27956
rect 11060 27940 11112 27946
rect 11060 27882 11112 27888
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 10980 25838 11008 26522
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10796 22234 10824 22510
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10612 22066 10732 22094
rect 10508 22034 10560 22040
rect 10704 21894 10732 22066
rect 10888 22030 10916 22510
rect 10980 22098 11008 25638
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10876 22024 10928 22030
rect 10928 21972 11008 21978
rect 10876 21966 11008 21972
rect 10888 21950 11008 21966
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10704 21622 10732 21830
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10520 20534 10548 20878
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10704 20346 10732 21286
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10796 20534 10824 20742
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10704 20318 10824 20346
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10704 19530 10732 19722
rect 10520 19502 10732 19530
rect 10414 17912 10470 17921
rect 10414 17847 10470 17856
rect 10428 17202 10456 17847
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10336 17054 10456 17082
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 9864 12378 9916 12384
rect 9968 12406 10180 12434
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 11762 9812 12174
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 9876 11354 9904 12378
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9508 9586 9536 9930
rect 9692 9586 9720 10066
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 9876 9160 9904 9386
rect 9324 9030 9444 9058
rect 9784 9132 9904 9160
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9232 6798 9260 8910
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9140 6616 9260 6644
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9232 3738 9260 6616
rect 9324 5914 9352 9030
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9416 7750 9444 8910
rect 9600 8634 9628 8910
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9784 8430 9812 9132
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9876 8838 9904 8978
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9862 8528 9918 8537
rect 9862 8463 9864 8472
rect 9916 8463 9918 8472
rect 9864 8434 9916 8440
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9416 6866 9444 7686
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9876 6866 9904 8298
rect 9968 7206 9996 12406
rect 10244 12306 10272 13874
rect 10336 13394 10364 16594
rect 10428 16182 10456 17054
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10428 15434 10456 15982
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10520 14600 10548 19502
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10428 14572 10548 14600
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10428 12434 10456 14572
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10336 12406 10456 12434
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10336 12102 10364 12406
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10060 11354 10088 11766
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10244 11218 10272 11766
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10336 10577 10364 12038
rect 10322 10568 10378 10577
rect 10322 10503 10378 10512
rect 10336 10266 10364 10503
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10048 9512 10100 9518
rect 10100 9472 10180 9500
rect 10048 9454 10100 9460
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 8838 10088 9318
rect 10152 9178 10180 9472
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10140 8968 10192 8974
rect 10138 8936 10140 8945
rect 10192 8936 10194 8945
rect 10138 8871 10194 8880
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10060 7342 10088 8774
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 6254 9904 6802
rect 9680 6248 9732 6254
rect 9678 6216 9680 6225
rect 9864 6248 9916 6254
rect 9732 6216 9734 6225
rect 9864 6190 9916 6196
rect 9678 6151 9734 6160
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9324 5642 9352 5850
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9416 4826 9444 5170
rect 9784 5114 9812 5714
rect 9876 5370 9904 6190
rect 9968 6186 9996 7142
rect 10060 6458 10088 7278
rect 10152 7002 10180 8871
rect 10244 8362 10272 10066
rect 10428 9874 10456 12310
rect 10336 9846 10456 9874
rect 10336 9217 10364 9846
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10428 9586 10456 9658
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10520 9330 10548 14418
rect 10612 12238 10640 19314
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 10704 17882 10732 19178
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17202 10732 17478
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10796 17082 10824 20318
rect 10888 20058 10916 21490
rect 10980 21350 11008 21950
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 11072 20369 11100 27882
rect 11532 27441 11560 27950
rect 11624 27946 11652 28999
rect 11612 27940 11664 27946
rect 11612 27882 11664 27888
rect 11612 27600 11664 27606
rect 11612 27542 11664 27548
rect 11518 27432 11574 27441
rect 11518 27367 11574 27376
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 11164 25265 11192 27270
rect 11230 27228 11538 27237
rect 11230 27226 11236 27228
rect 11292 27226 11316 27228
rect 11372 27226 11396 27228
rect 11452 27226 11476 27228
rect 11532 27226 11538 27228
rect 11292 27174 11294 27226
rect 11474 27174 11476 27226
rect 11230 27172 11236 27174
rect 11292 27172 11316 27174
rect 11372 27172 11396 27174
rect 11452 27172 11476 27174
rect 11532 27172 11538 27174
rect 11230 27163 11538 27172
rect 11428 26988 11480 26994
rect 11428 26930 11480 26936
rect 11440 26586 11468 26930
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11532 26586 11560 26726
rect 11428 26580 11480 26586
rect 11428 26522 11480 26528
rect 11520 26580 11572 26586
rect 11520 26522 11572 26528
rect 11230 26140 11538 26149
rect 11230 26138 11236 26140
rect 11292 26138 11316 26140
rect 11372 26138 11396 26140
rect 11452 26138 11476 26140
rect 11532 26138 11538 26140
rect 11292 26086 11294 26138
rect 11474 26086 11476 26138
rect 11230 26084 11236 26086
rect 11292 26084 11316 26086
rect 11372 26084 11396 26086
rect 11452 26084 11476 26086
rect 11532 26084 11538 26086
rect 11230 26075 11538 26084
rect 11150 25256 11206 25265
rect 11150 25191 11206 25200
rect 11230 25052 11538 25061
rect 11230 25050 11236 25052
rect 11292 25050 11316 25052
rect 11372 25050 11396 25052
rect 11452 25050 11476 25052
rect 11532 25050 11538 25052
rect 11292 24998 11294 25050
rect 11474 24998 11476 25050
rect 11230 24996 11236 24998
rect 11292 24996 11316 24998
rect 11372 24996 11396 24998
rect 11452 24996 11476 24998
rect 11532 24996 11538 24998
rect 11230 24987 11538 24996
rect 11244 24948 11296 24954
rect 11244 24890 11296 24896
rect 11256 24410 11284 24890
rect 11624 24698 11652 27542
rect 11716 27538 11744 32932
rect 11888 32836 11940 32842
rect 11888 32778 11940 32784
rect 11900 31482 11928 32778
rect 11992 32774 12020 34614
rect 12084 33946 12112 34904
rect 12348 34886 12400 34892
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12440 34604 12492 34610
rect 12440 34546 12492 34552
rect 12268 34513 12296 34546
rect 12348 34536 12400 34542
rect 12254 34504 12310 34513
rect 12348 34478 12400 34484
rect 12254 34439 12310 34448
rect 12084 33918 12204 33946
rect 12072 33856 12124 33862
rect 12072 33798 12124 33804
rect 11980 32768 12032 32774
rect 11980 32710 12032 32716
rect 11980 32496 12032 32502
rect 11980 32438 12032 32444
rect 11992 31958 12020 32438
rect 11980 31952 12032 31958
rect 11980 31894 12032 31900
rect 11980 31816 12032 31822
rect 11978 31784 11980 31793
rect 12032 31784 12034 31793
rect 11978 31719 12034 31728
rect 11888 31476 11940 31482
rect 11888 31418 11940 31424
rect 11886 31376 11942 31385
rect 11886 31311 11888 31320
rect 11940 31311 11942 31320
rect 11888 31282 11940 31288
rect 12084 31260 12112 33798
rect 12176 33658 12204 33918
rect 12164 33652 12216 33658
rect 12164 33594 12216 33600
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 12176 33425 12204 33458
rect 12162 33416 12218 33425
rect 12162 33351 12218 33360
rect 12164 32768 12216 32774
rect 12164 32710 12216 32716
rect 12176 31362 12204 32710
rect 12360 32473 12388 34478
rect 12452 33114 12480 34546
rect 12440 33108 12492 33114
rect 12440 33050 12492 33056
rect 12440 32836 12492 32842
rect 12440 32778 12492 32784
rect 12346 32464 12402 32473
rect 12346 32399 12402 32408
rect 12348 32020 12400 32026
rect 12452 32008 12480 32778
rect 12544 32450 12572 34886
rect 12636 32609 12664 36230
rect 13266 36207 13322 36216
rect 12716 36100 12768 36106
rect 12716 36042 12768 36048
rect 12992 36100 13044 36106
rect 12992 36042 13044 36048
rect 13176 36100 13228 36106
rect 13176 36042 13228 36048
rect 12728 35170 12756 36042
rect 13004 35578 13032 36042
rect 13188 35630 13216 36042
rect 13268 36032 13320 36038
rect 13268 35974 13320 35980
rect 13280 35737 13308 35974
rect 13266 35728 13322 35737
rect 13266 35663 13322 35672
rect 12820 35550 13032 35578
rect 13176 35624 13228 35630
rect 13176 35566 13228 35572
rect 12820 35290 12848 35550
rect 12944 35388 13252 35397
rect 12944 35386 12950 35388
rect 13006 35386 13030 35388
rect 13086 35386 13110 35388
rect 13166 35386 13190 35388
rect 13246 35386 13252 35388
rect 13006 35334 13008 35386
rect 13188 35334 13190 35386
rect 12944 35332 12950 35334
rect 13006 35332 13030 35334
rect 13086 35332 13110 35334
rect 13166 35332 13190 35334
rect 13246 35332 13252 35334
rect 12944 35323 13252 35332
rect 12808 35284 12860 35290
rect 12808 35226 12860 35232
rect 12728 35142 12848 35170
rect 12820 33998 12848 35142
rect 13268 34944 13320 34950
rect 13268 34886 13320 34892
rect 12944 34300 13252 34309
rect 12944 34298 12950 34300
rect 13006 34298 13030 34300
rect 13086 34298 13110 34300
rect 13166 34298 13190 34300
rect 13246 34298 13252 34300
rect 13006 34246 13008 34298
rect 13188 34246 13190 34298
rect 12944 34244 12950 34246
rect 13006 34244 13030 34246
rect 13086 34244 13110 34246
rect 13166 34244 13190 34246
rect 13246 34244 13252 34246
rect 12944 34235 13252 34244
rect 13280 34105 13308 34886
rect 13360 34604 13412 34610
rect 13360 34546 13412 34552
rect 13266 34096 13322 34105
rect 13266 34031 13322 34040
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12992 33992 13044 33998
rect 12992 33934 13044 33940
rect 12716 33924 12768 33930
rect 12716 33866 12768 33872
rect 12728 32842 12756 33866
rect 13004 33318 13032 33934
rect 13268 33856 13320 33862
rect 13268 33798 13320 33804
rect 12900 33312 12952 33318
rect 12820 33272 12900 33300
rect 12716 32836 12768 32842
rect 12716 32778 12768 32784
rect 12622 32600 12678 32609
rect 12622 32535 12678 32544
rect 12544 32422 12756 32450
rect 12532 32224 12584 32230
rect 12532 32166 12584 32172
rect 12624 32224 12676 32230
rect 12624 32166 12676 32172
rect 12400 31980 12480 32008
rect 12348 31962 12400 31968
rect 12544 31958 12572 32166
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12360 31385 12388 31758
rect 12346 31376 12402 31385
rect 12176 31334 12296 31362
rect 12164 31272 12216 31278
rect 12084 31232 12164 31260
rect 12164 31214 12216 31220
rect 11888 31204 11940 31210
rect 11888 31146 11940 31152
rect 11796 30796 11848 30802
rect 11796 30738 11848 30744
rect 11808 29753 11836 30738
rect 11794 29744 11850 29753
rect 11794 29679 11850 29688
rect 11900 28506 11928 31146
rect 12162 30832 12218 30841
rect 12268 30818 12296 31334
rect 12346 31311 12402 31320
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12532 31272 12584 31278
rect 12532 31214 12584 31220
rect 12636 31226 12664 32166
rect 12728 31346 12756 32422
rect 12820 31906 12848 33272
rect 12900 33254 12952 33260
rect 12992 33312 13044 33318
rect 12992 33254 13044 33260
rect 12944 33212 13252 33221
rect 12944 33210 12950 33212
rect 13006 33210 13030 33212
rect 13086 33210 13110 33212
rect 13166 33210 13190 33212
rect 13246 33210 13252 33212
rect 13006 33158 13008 33210
rect 13188 33158 13190 33210
rect 12944 33156 12950 33158
rect 13006 33156 13030 33158
rect 13086 33156 13110 33158
rect 13166 33156 13190 33158
rect 13246 33156 13252 33158
rect 12944 33147 13252 33156
rect 12992 32768 13044 32774
rect 12992 32710 13044 32716
rect 13004 32570 13032 32710
rect 12992 32564 13044 32570
rect 12992 32506 13044 32512
rect 12992 32428 13044 32434
rect 12992 32370 13044 32376
rect 13004 32337 13032 32370
rect 12990 32328 13046 32337
rect 12990 32263 13046 32272
rect 12944 32124 13252 32133
rect 12944 32122 12950 32124
rect 13006 32122 13030 32124
rect 13086 32122 13110 32124
rect 13166 32122 13190 32124
rect 13246 32122 13252 32124
rect 13006 32070 13008 32122
rect 13188 32070 13190 32122
rect 12944 32068 12950 32070
rect 13006 32068 13030 32070
rect 13086 32068 13110 32070
rect 13166 32068 13190 32070
rect 13246 32068 13252 32070
rect 12944 32059 13252 32068
rect 12820 31878 13216 31906
rect 13188 31822 13216 31878
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 13084 31816 13136 31822
rect 13084 31758 13136 31764
rect 13176 31816 13228 31822
rect 13176 31758 13228 31764
rect 12716 31340 12768 31346
rect 12716 31282 12768 31288
rect 12218 30790 12296 30818
rect 12162 30767 12218 30776
rect 12452 30784 12480 31214
rect 12544 31142 12572 31214
rect 12636 31198 12756 31226
rect 12532 31136 12584 31142
rect 12532 31078 12584 31084
rect 12728 30870 12756 31198
rect 12912 31192 12940 31758
rect 12820 31164 12940 31192
rect 12716 30864 12768 30870
rect 12716 30806 12768 30812
rect 12820 30802 12848 31164
rect 13096 31124 13124 31758
rect 13280 31278 13308 33798
rect 13372 33153 13400 34546
rect 13464 34490 13492 36502
rect 13648 35850 13676 36790
rect 13726 36751 13782 36760
rect 13820 36780 13872 36786
rect 13820 36722 13872 36728
rect 14004 36780 14056 36786
rect 14004 36722 14056 36728
rect 13728 36576 13780 36582
rect 13728 36518 13780 36524
rect 13740 36145 13768 36518
rect 13832 36281 13860 36722
rect 13818 36272 13874 36281
rect 13818 36207 13874 36216
rect 13726 36136 13782 36145
rect 13726 36071 13782 36080
rect 13648 35822 13768 35850
rect 13544 35692 13596 35698
rect 13544 35634 13596 35640
rect 13636 35692 13688 35698
rect 13636 35634 13688 35640
rect 13556 34746 13584 35634
rect 13648 35057 13676 35634
rect 13634 35048 13690 35057
rect 13634 34983 13690 34992
rect 13544 34740 13596 34746
rect 13544 34682 13596 34688
rect 13542 34640 13598 34649
rect 13542 34575 13544 34584
rect 13596 34575 13598 34584
rect 13544 34546 13596 34552
rect 13464 34462 13676 34490
rect 13544 33856 13596 33862
rect 13544 33798 13596 33804
rect 13358 33144 13414 33153
rect 13358 33079 13414 33088
rect 13360 32836 13412 32842
rect 13360 32778 13412 32784
rect 13268 31272 13320 31278
rect 13372 31249 13400 32778
rect 13556 32570 13584 33798
rect 13648 33697 13676 34462
rect 13634 33688 13690 33697
rect 13634 33623 13690 33632
rect 13740 33538 13768 35822
rect 13820 35488 13872 35494
rect 13820 35430 13872 35436
rect 13832 34649 13860 35430
rect 13818 34640 13874 34649
rect 13818 34575 13874 34584
rect 13820 34400 13872 34406
rect 13820 34342 13872 34348
rect 13648 33510 13768 33538
rect 13648 33017 13676 33510
rect 13832 33289 13860 34342
rect 14016 33522 14044 36722
rect 14188 36168 14240 36174
rect 14188 36110 14240 36116
rect 14200 35834 14228 36110
rect 14188 35828 14240 35834
rect 14188 35770 14240 35776
rect 14292 35034 14320 41386
rect 15028 41386 15148 41414
rect 14657 41372 14965 41381
rect 14657 41370 14663 41372
rect 14719 41370 14743 41372
rect 14799 41370 14823 41372
rect 14879 41370 14903 41372
rect 14959 41370 14965 41372
rect 14719 41318 14721 41370
rect 14901 41318 14903 41370
rect 14657 41316 14663 41318
rect 14719 41316 14743 41318
rect 14799 41316 14823 41318
rect 14879 41316 14903 41318
rect 14959 41316 14965 41318
rect 14657 41307 14965 41316
rect 14657 40284 14965 40293
rect 14657 40282 14663 40284
rect 14719 40282 14743 40284
rect 14799 40282 14823 40284
rect 14879 40282 14903 40284
rect 14959 40282 14965 40284
rect 14719 40230 14721 40282
rect 14901 40230 14903 40282
rect 14657 40228 14663 40230
rect 14719 40228 14743 40230
rect 14799 40228 14823 40230
rect 14879 40228 14903 40230
rect 14959 40228 14965 40230
rect 14657 40219 14965 40228
rect 14372 39296 14424 39302
rect 14372 39238 14424 39244
rect 14384 38729 14412 39238
rect 14657 39196 14965 39205
rect 14657 39194 14663 39196
rect 14719 39194 14743 39196
rect 14799 39194 14823 39196
rect 14879 39194 14903 39196
rect 14959 39194 14965 39196
rect 14719 39142 14721 39194
rect 14901 39142 14903 39194
rect 14657 39140 14663 39142
rect 14719 39140 14743 39142
rect 14799 39140 14823 39142
rect 14879 39140 14903 39142
rect 14959 39140 14965 39142
rect 14657 39131 14965 39140
rect 14370 38720 14426 38729
rect 14370 38655 14426 38664
rect 14372 38208 14424 38214
rect 14372 38150 14424 38156
rect 14384 37641 14412 38150
rect 14657 38108 14965 38117
rect 14657 38106 14663 38108
rect 14719 38106 14743 38108
rect 14799 38106 14823 38108
rect 14879 38106 14903 38108
rect 14959 38106 14965 38108
rect 14719 38054 14721 38106
rect 14901 38054 14903 38106
rect 14657 38052 14663 38054
rect 14719 38052 14743 38054
rect 14799 38052 14823 38054
rect 14879 38052 14903 38054
rect 14959 38052 14965 38054
rect 14657 38043 14965 38052
rect 14370 37632 14426 37641
rect 14370 37567 14426 37576
rect 14372 37120 14424 37126
rect 14372 37062 14424 37068
rect 14384 36553 14412 37062
rect 14657 37020 14965 37029
rect 14657 37018 14663 37020
rect 14719 37018 14743 37020
rect 14799 37018 14823 37020
rect 14879 37018 14903 37020
rect 14959 37018 14965 37020
rect 14719 36966 14721 37018
rect 14901 36966 14903 37018
rect 14657 36964 14663 36966
rect 14719 36964 14743 36966
rect 14799 36964 14823 36966
rect 14879 36964 14903 36966
rect 14959 36964 14965 36966
rect 14657 36955 14965 36964
rect 14370 36544 14426 36553
rect 14370 36479 14426 36488
rect 14657 35932 14965 35941
rect 14657 35930 14663 35932
rect 14719 35930 14743 35932
rect 14799 35930 14823 35932
rect 14879 35930 14903 35932
rect 14959 35930 14965 35932
rect 14719 35878 14721 35930
rect 14901 35878 14903 35930
rect 14657 35876 14663 35878
rect 14719 35876 14743 35878
rect 14799 35876 14823 35878
rect 14879 35876 14903 35878
rect 14959 35876 14965 35878
rect 14657 35867 14965 35876
rect 14464 35624 14516 35630
rect 14464 35566 14516 35572
rect 14476 35193 14504 35566
rect 14462 35184 14518 35193
rect 14462 35119 14518 35128
rect 14292 35006 14504 35034
rect 14096 34604 14148 34610
rect 14096 34546 14148 34552
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 14108 33402 14136 34546
rect 14280 33992 14332 33998
rect 14280 33934 14332 33940
rect 13924 33374 14136 33402
rect 13818 33280 13874 33289
rect 13818 33215 13874 33224
rect 13728 33040 13780 33046
rect 13634 33008 13690 33017
rect 13728 32982 13780 32988
rect 13634 32943 13690 32952
rect 13544 32564 13596 32570
rect 13544 32506 13596 32512
rect 13544 32224 13596 32230
rect 13544 32166 13596 32172
rect 13452 31680 13504 31686
rect 13452 31622 13504 31628
rect 13464 31414 13492 31622
rect 13452 31408 13504 31414
rect 13452 31350 13504 31356
rect 13268 31214 13320 31220
rect 13358 31240 13414 31249
rect 13358 31175 13414 31184
rect 13096 31096 13492 31124
rect 12944 31036 13252 31045
rect 12944 31034 12950 31036
rect 13006 31034 13030 31036
rect 13086 31034 13110 31036
rect 13166 31034 13190 31036
rect 13246 31034 13252 31036
rect 13006 30982 13008 31034
rect 13188 30982 13190 31034
rect 12944 30980 12950 30982
rect 13006 30980 13030 30982
rect 13086 30980 13110 30982
rect 13166 30980 13190 30982
rect 13246 30980 13252 30982
rect 12944 30971 13252 30980
rect 12624 30796 12676 30802
rect 12452 30756 12624 30784
rect 11980 30660 12032 30666
rect 11980 30602 12032 30608
rect 11808 28478 11928 28506
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 11716 27130 11744 27270
rect 11704 27124 11756 27130
rect 11704 27066 11756 27072
rect 11704 26920 11756 26926
rect 11704 26862 11756 26868
rect 11348 24670 11652 24698
rect 11244 24404 11296 24410
rect 11244 24346 11296 24352
rect 11348 24052 11376 24670
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11440 24342 11468 24550
rect 11428 24336 11480 24342
rect 11428 24278 11480 24284
rect 11532 24120 11560 24550
rect 11532 24092 11652 24120
rect 11164 24024 11376 24052
rect 11164 23118 11192 24024
rect 11230 23964 11538 23973
rect 11230 23962 11236 23964
rect 11292 23962 11316 23964
rect 11372 23962 11396 23964
rect 11452 23962 11476 23964
rect 11532 23962 11538 23964
rect 11292 23910 11294 23962
rect 11474 23910 11476 23962
rect 11230 23908 11236 23910
rect 11292 23908 11316 23910
rect 11372 23908 11396 23910
rect 11452 23908 11476 23910
rect 11532 23908 11538 23910
rect 11230 23899 11538 23908
rect 11624 23202 11652 24092
rect 11716 24070 11744 26862
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11624 23186 11744 23202
rect 11624 23180 11756 23186
rect 11624 23174 11704 23180
rect 11704 23122 11756 23128
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11164 22681 11192 23054
rect 11230 22876 11538 22885
rect 11230 22874 11236 22876
rect 11292 22874 11316 22876
rect 11372 22874 11396 22876
rect 11452 22874 11476 22876
rect 11532 22874 11538 22876
rect 11292 22822 11294 22874
rect 11474 22822 11476 22874
rect 11230 22820 11236 22822
rect 11292 22820 11316 22822
rect 11372 22820 11396 22822
rect 11452 22820 11476 22822
rect 11532 22820 11538 22822
rect 11230 22811 11538 22820
rect 11150 22672 11206 22681
rect 11150 22607 11206 22616
rect 11808 22094 11836 28478
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11900 26489 11928 28358
rect 11992 27577 12020 30602
rect 12072 30592 12124 30598
rect 12072 30534 12124 30540
rect 12440 30592 12492 30598
rect 12440 30534 12492 30540
rect 12084 28994 12112 30534
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12268 30161 12296 30194
rect 12254 30152 12310 30161
rect 12254 30087 12310 30096
rect 12164 30048 12216 30054
rect 12164 29990 12216 29996
rect 12176 29170 12204 29990
rect 12346 29880 12402 29889
rect 12346 29815 12402 29824
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12268 29209 12296 29242
rect 12254 29200 12310 29209
rect 12162 29164 12214 29170
rect 12254 29135 12310 29144
rect 12162 29106 12214 29112
rect 12084 28966 12204 28994
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 12084 27674 12112 28494
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 11978 27568 12034 27577
rect 12176 27538 12204 28966
rect 12256 28960 12308 28966
rect 12256 28902 12308 28908
rect 12268 28218 12296 28902
rect 12256 28212 12308 28218
rect 12256 28154 12308 28160
rect 12360 28121 12388 29815
rect 12346 28112 12402 28121
rect 12346 28047 12402 28056
rect 12452 27690 12480 30534
rect 12544 27878 12572 30756
rect 12624 30738 12676 30744
rect 12808 30796 12860 30802
rect 12808 30738 12860 30744
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 13188 30138 13216 30670
rect 13188 30110 13308 30138
rect 12624 30048 12676 30054
rect 12900 30048 12952 30054
rect 12624 29990 12676 29996
rect 12820 30008 12900 30036
rect 12636 29850 12664 29990
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12624 29708 12676 29714
rect 12624 29650 12676 29656
rect 12636 29617 12664 29650
rect 12622 29608 12678 29617
rect 12622 29543 12678 29552
rect 12624 29504 12676 29510
rect 12624 29446 12676 29452
rect 12636 29306 12664 29446
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 12622 29064 12678 29073
rect 12622 28999 12678 29008
rect 12636 28694 12664 28999
rect 12716 28960 12768 28966
rect 12716 28902 12768 28908
rect 12624 28688 12676 28694
rect 12624 28630 12676 28636
rect 12728 28540 12756 28902
rect 12820 28694 12848 30008
rect 12900 29990 12952 29996
rect 12944 29948 13252 29957
rect 12944 29946 12950 29948
rect 13006 29946 13030 29948
rect 13086 29946 13110 29948
rect 13166 29946 13190 29948
rect 13246 29946 13252 29948
rect 13006 29894 13008 29946
rect 13188 29894 13190 29946
rect 12944 29892 12950 29894
rect 13006 29892 13030 29894
rect 13086 29892 13110 29894
rect 13166 29892 13190 29894
rect 13246 29892 13252 29894
rect 12944 29883 13252 29892
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 13004 29102 13032 29514
rect 12992 29096 13044 29102
rect 13176 29096 13228 29102
rect 12992 29038 13044 29044
rect 13174 29064 13176 29073
rect 13228 29064 13230 29073
rect 13174 28999 13230 29008
rect 12944 28860 13252 28869
rect 12944 28858 12950 28860
rect 13006 28858 13030 28860
rect 13086 28858 13110 28860
rect 13166 28858 13190 28860
rect 13246 28858 13252 28860
rect 13006 28806 13008 28858
rect 13188 28806 13190 28858
rect 12944 28804 12950 28806
rect 13006 28804 13030 28806
rect 13086 28804 13110 28806
rect 13166 28804 13190 28806
rect 13246 28804 13252 28806
rect 12944 28795 13252 28804
rect 12808 28688 12860 28694
rect 12808 28630 12860 28636
rect 13176 28620 13228 28626
rect 13176 28562 13228 28568
rect 12992 28552 13044 28558
rect 12636 28512 12992 28540
rect 12532 27872 12584 27878
rect 12532 27814 12584 27820
rect 12452 27662 12572 27690
rect 11978 27503 12034 27512
rect 12164 27532 12216 27538
rect 12164 27474 12216 27480
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 12452 27441 12480 27474
rect 12438 27432 12494 27441
rect 12360 27390 12438 27418
rect 12072 26512 12124 26518
rect 11886 26480 11942 26489
rect 12072 26454 12124 26460
rect 11886 26415 11942 26424
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11900 24857 11928 25638
rect 11980 25220 12032 25226
rect 11980 25162 12032 25168
rect 11886 24848 11942 24857
rect 11886 24783 11942 24792
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 11900 24274 11928 24346
rect 11992 24313 12020 25162
rect 12084 24954 12112 26454
rect 12164 26376 12216 26382
rect 12216 26336 12296 26364
rect 12164 26318 12216 26324
rect 12164 25832 12216 25838
rect 12268 25809 12296 26336
rect 12164 25774 12216 25780
rect 12254 25800 12310 25809
rect 12072 24948 12124 24954
rect 12072 24890 12124 24896
rect 12176 24410 12204 25774
rect 12254 25735 12310 25744
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 11978 24304 12034 24313
rect 11888 24268 11940 24274
rect 11978 24239 12034 24248
rect 11888 24210 11940 24216
rect 11900 22234 11928 24210
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 11980 23180 12032 23186
rect 11980 23122 12032 23128
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11808 22066 11928 22094
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11230 21788 11538 21797
rect 11230 21786 11236 21788
rect 11292 21786 11316 21788
rect 11372 21786 11396 21788
rect 11452 21786 11476 21788
rect 11532 21786 11538 21788
rect 11292 21734 11294 21786
rect 11474 21734 11476 21786
rect 11230 21732 11236 21734
rect 11292 21732 11316 21734
rect 11372 21732 11396 21734
rect 11452 21732 11476 21734
rect 11532 21732 11538 21734
rect 11230 21723 11538 21732
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11164 20602 11192 20742
rect 11230 20700 11538 20709
rect 11230 20698 11236 20700
rect 11292 20698 11316 20700
rect 11372 20698 11396 20700
rect 11452 20698 11476 20700
rect 11532 20698 11538 20700
rect 11292 20646 11294 20698
rect 11474 20646 11476 20698
rect 11230 20644 11236 20646
rect 11292 20644 11316 20646
rect 11372 20644 11396 20646
rect 11452 20644 11476 20646
rect 11532 20644 11538 20646
rect 11230 20635 11538 20644
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11624 20534 11652 21830
rect 11794 21448 11850 21457
rect 11794 21383 11850 21392
rect 11612 20528 11664 20534
rect 11612 20470 11664 20476
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11058 20360 11114 20369
rect 11058 20295 11114 20304
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10888 19378 10916 19450
rect 10966 19408 11022 19417
rect 10876 19372 10928 19378
rect 10966 19343 11022 19352
rect 10876 19314 10928 19320
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 18426 10916 18566
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10888 17542 10916 17750
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10876 17128 10928 17134
rect 10796 17076 10876 17082
rect 10796 17070 10928 17076
rect 10796 17054 10916 17070
rect 10796 16114 10824 17054
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16658 10916 16934
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 14482 10732 15302
rect 10796 14958 10824 15370
rect 10888 15008 10916 16594
rect 10980 15416 11008 19343
rect 11072 16572 11100 20198
rect 11164 19514 11192 20402
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11336 20324 11388 20330
rect 11336 20266 11388 20272
rect 11348 19922 11376 20266
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11230 19612 11538 19621
rect 11230 19610 11236 19612
rect 11292 19610 11316 19612
rect 11372 19610 11396 19612
rect 11452 19610 11476 19612
rect 11532 19610 11538 19612
rect 11292 19558 11294 19610
rect 11474 19558 11476 19610
rect 11230 19556 11236 19558
rect 11292 19556 11316 19558
rect 11372 19556 11396 19558
rect 11452 19556 11476 19558
rect 11532 19556 11538 19558
rect 11230 19547 11538 19556
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 11624 18834 11652 20334
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11716 19310 11744 20198
rect 11808 20058 11836 21383
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18834 11744 19110
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11794 18728 11850 18737
rect 11612 18692 11664 18698
rect 11612 18634 11664 18640
rect 11716 18686 11794 18714
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 18426 11192 18566
rect 11230 18524 11538 18533
rect 11230 18522 11236 18524
rect 11292 18522 11316 18524
rect 11372 18522 11396 18524
rect 11452 18522 11476 18524
rect 11532 18522 11538 18524
rect 11292 18470 11294 18522
rect 11474 18470 11476 18522
rect 11230 18468 11236 18470
rect 11292 18468 11316 18470
rect 11372 18468 11396 18470
rect 11452 18468 11476 18470
rect 11532 18468 11538 18470
rect 11230 18459 11538 18468
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11164 17785 11192 18226
rect 11426 18184 11482 18193
rect 11426 18119 11482 18128
rect 11150 17776 11206 17785
rect 11150 17711 11206 17720
rect 11440 17678 11468 18119
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11532 17524 11560 17614
rect 11164 17496 11560 17524
rect 11164 17116 11192 17496
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11244 17128 11296 17134
rect 11164 17088 11244 17116
rect 11440 17105 11468 17206
rect 11244 17070 11296 17076
rect 11426 17096 11482 17105
rect 11152 16584 11204 16590
rect 11072 16544 11152 16572
rect 11152 16526 11204 16532
rect 11256 16436 11284 17070
rect 11426 17031 11482 17040
rect 11164 16408 11284 16436
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 15706 11100 16050
rect 11164 16046 11192 16408
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15706 11192 15846
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11532 15450 11560 15982
rect 11624 15910 11652 18634
rect 11716 17882 11744 18686
rect 11900 18714 11928 22066
rect 11992 22030 12020 23122
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11992 21010 12020 21966
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 11978 20904 12034 20913
rect 11978 20839 12034 20848
rect 11992 18970 12020 20839
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11900 18686 12020 18714
rect 11794 18663 11850 18672
rect 11888 18624 11940 18630
rect 11794 18592 11850 18601
rect 11888 18566 11940 18572
rect 11794 18527 11850 18536
rect 11808 18034 11836 18527
rect 11900 18426 11928 18566
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11808 18006 11928 18034
rect 11794 17912 11850 17921
rect 11704 17876 11756 17882
rect 11794 17847 11850 17856
rect 11704 17818 11756 17824
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17241 11744 17682
rect 11808 17513 11836 17847
rect 11794 17504 11850 17513
rect 11794 17439 11850 17448
rect 11702 17232 11758 17241
rect 11702 17167 11758 17176
rect 11794 17096 11850 17105
rect 11794 17031 11850 17040
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11716 16658 11744 16934
rect 11808 16794 11836 17031
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11532 15422 11744 15450
rect 10980 15388 11100 15416
rect 10888 14980 11008 15008
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14618 10824 14758
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10704 12442 10732 13670
rect 10796 13138 10824 14350
rect 10796 13110 10916 13138
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10612 11014 10640 12174
rect 10704 11762 10732 12242
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10796 10962 10824 12786
rect 10888 11354 10916 13110
rect 10980 12374 11008 14980
rect 11072 14521 11100 15388
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11058 14512 11114 14521
rect 11058 14447 11114 14456
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 11072 12850 11100 13942
rect 11164 13410 11192 14418
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 14278 11376 14350
rect 11336 14272 11388 14278
rect 11532 14260 11560 14554
rect 11624 14482 11652 15302
rect 11716 14498 11744 15422
rect 11808 14618 11836 16594
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11612 14476 11664 14482
rect 11716 14470 11836 14498
rect 11612 14418 11664 14424
rect 11808 14328 11836 14470
rect 11714 14300 11836 14328
rect 11714 14260 11742 14300
rect 11532 14232 11652 14260
rect 11714 14232 11744 14260
rect 11336 14214 11388 14220
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 11164 13382 11284 13410
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 11164 11694 11192 13262
rect 11256 13190 11284 13382
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11164 11506 11192 11630
rect 11164 11478 11284 11506
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11256 11286 11284 11478
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10612 10130 10640 10950
rect 10796 10934 10916 10962
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10612 10033 10640 10066
rect 10598 10024 10654 10033
rect 10598 9959 10654 9968
rect 10612 9586 10640 9959
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10428 9302 10548 9330
rect 10322 9208 10378 9217
rect 10322 9143 10378 9152
rect 10336 9042 10364 9143
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10152 6866 10180 6938
rect 10336 6866 10364 8978
rect 10428 7342 10456 9302
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10520 8498 10548 9114
rect 10704 8498 10732 10474
rect 10796 10062 10824 10746
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10796 9722 10824 9998
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10888 9602 10916 10934
rect 11072 10713 11100 11086
rect 11058 10704 11114 10713
rect 11058 10639 11114 10648
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9722 11008 9862
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10796 9574 10916 9602
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 7698 10732 8434
rect 10612 7670 10732 7698
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10428 6254 10456 7278
rect 10612 6866 10640 7670
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10704 7410 10732 7482
rect 10796 7426 10824 9574
rect 10876 9512 10928 9518
rect 10928 9472 11008 9500
rect 10876 9454 10928 9460
rect 10874 9072 10930 9081
rect 10980 9042 11008 9472
rect 11072 9178 11100 10202
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10874 9007 10930 9016
rect 10968 9036 11020 9042
rect 10888 8294 10916 9007
rect 10968 8978 11020 8984
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 7886 10916 8230
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10980 7546 11008 8978
rect 11164 8945 11192 11222
rect 11624 11082 11652 14232
rect 11716 14006 11744 14232
rect 11794 14240 11850 14249
rect 11794 14175 11850 14184
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11808 13938 11836 14175
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11702 13832 11758 13841
rect 11702 13767 11758 13776
rect 11716 12986 11744 13767
rect 11900 13394 11928 18006
rect 11992 16658 12020 18686
rect 12084 17746 12112 23598
rect 12176 22137 12204 23666
rect 12268 23662 12296 25735
rect 12360 25498 12388 27390
rect 12438 27367 12494 27376
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12452 26518 12480 26930
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12452 25838 12480 26318
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12348 25492 12400 25498
rect 12348 25434 12400 25440
rect 12544 25378 12572 27662
rect 12636 26450 12664 28512
rect 12992 28494 13044 28500
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12728 27441 12756 28018
rect 13188 27878 13216 28562
rect 12808 27872 12860 27878
rect 12808 27814 12860 27820
rect 13176 27872 13228 27878
rect 13176 27814 13228 27820
rect 12714 27432 12770 27441
rect 12714 27367 12770 27376
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12728 26790 12756 26930
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12820 26518 12848 27814
rect 12944 27772 13252 27781
rect 12944 27770 12950 27772
rect 13006 27770 13030 27772
rect 13086 27770 13110 27772
rect 13166 27770 13190 27772
rect 13246 27770 13252 27772
rect 13006 27718 13008 27770
rect 13188 27718 13190 27770
rect 12944 27716 12950 27718
rect 13006 27716 13030 27718
rect 13086 27716 13110 27718
rect 13166 27716 13190 27718
rect 13246 27716 13252 27718
rect 12944 27707 13252 27716
rect 13280 27418 13308 30110
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13188 27390 13308 27418
rect 13188 26858 13216 27390
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13176 26852 13228 26858
rect 13176 26794 13228 26800
rect 12944 26684 13252 26693
rect 12944 26682 12950 26684
rect 13006 26682 13030 26684
rect 13086 26682 13110 26684
rect 13166 26682 13190 26684
rect 13246 26682 13252 26684
rect 13006 26630 13008 26682
rect 13188 26630 13190 26682
rect 12944 26628 12950 26630
rect 13006 26628 13030 26630
rect 13086 26628 13110 26630
rect 13166 26628 13190 26630
rect 13246 26628 13252 26630
rect 12944 26619 13252 26628
rect 13280 26586 13308 27270
rect 13372 27062 13400 28358
rect 13464 27606 13492 31096
rect 13556 30569 13584 32166
rect 13636 31272 13688 31278
rect 13636 31214 13688 31220
rect 13648 30802 13676 31214
rect 13636 30796 13688 30802
rect 13636 30738 13688 30744
rect 13542 30560 13598 30569
rect 13542 30495 13598 30504
rect 13544 29776 13596 29782
rect 13544 29718 13596 29724
rect 13556 29578 13584 29718
rect 13740 29646 13768 32982
rect 13818 31920 13874 31929
rect 13818 31855 13820 31864
rect 13872 31855 13874 31864
rect 13820 31826 13872 31832
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13544 29572 13596 29578
rect 13544 29514 13596 29520
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13544 28960 13596 28966
rect 13544 28902 13596 28908
rect 13556 28082 13584 28902
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13648 27985 13676 29446
rect 13832 29209 13860 31078
rect 13924 30938 13952 33374
rect 14004 33312 14056 33318
rect 14004 33254 14056 33260
rect 14188 33312 14240 33318
rect 14188 33254 14240 33260
rect 14016 32337 14044 33254
rect 14200 32745 14228 33254
rect 14292 33046 14320 33934
rect 14280 33040 14332 33046
rect 14280 32982 14332 32988
rect 14280 32904 14332 32910
rect 14280 32846 14332 32852
rect 14186 32736 14242 32745
rect 14186 32671 14242 32680
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14002 32328 14058 32337
rect 14002 32263 14058 32272
rect 14004 32224 14056 32230
rect 14004 32166 14056 32172
rect 14016 31958 14044 32166
rect 14004 31952 14056 31958
rect 14004 31894 14056 31900
rect 14108 31754 14136 32370
rect 14188 32360 14240 32366
rect 14188 32302 14240 32308
rect 14016 31726 14136 31754
rect 13912 30932 13964 30938
rect 13912 30874 13964 30880
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 13818 29200 13874 29209
rect 13818 29135 13874 29144
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13634 27976 13690 27985
rect 13634 27911 13690 27920
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13452 27600 13504 27606
rect 13452 27542 13504 27548
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13360 27056 13412 27062
rect 13360 26998 13412 27004
rect 13360 26852 13412 26858
rect 13360 26794 13412 26800
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 12808 26512 12860 26518
rect 13372 26466 13400 26794
rect 12808 26454 12860 26460
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 13096 26438 13400 26466
rect 12452 25350 12572 25378
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 12162 22128 12218 22137
rect 12162 22063 12218 22072
rect 12452 21894 12480 25350
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12544 24410 12572 24550
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12636 24274 12664 26386
rect 12992 25900 13044 25906
rect 13096 25888 13124 26438
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13044 25860 13124 25888
rect 12992 25842 13044 25848
rect 13188 25838 13216 26318
rect 13360 26036 13412 26042
rect 13360 25978 13412 25984
rect 13176 25832 13228 25838
rect 13176 25774 13228 25780
rect 12808 25764 12860 25770
rect 12808 25706 12860 25712
rect 13268 25764 13320 25770
rect 13268 25706 13320 25712
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12176 21049 12204 21490
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12268 21185 12296 21422
rect 12452 21350 12480 21626
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12254 21176 12310 21185
rect 12544 21162 12572 23734
rect 12820 23662 12848 25706
rect 12944 25596 13252 25605
rect 12944 25594 12950 25596
rect 13006 25594 13030 25596
rect 13086 25594 13110 25596
rect 13166 25594 13190 25596
rect 13246 25594 13252 25596
rect 13006 25542 13008 25594
rect 13188 25542 13190 25594
rect 12944 25540 12950 25542
rect 13006 25540 13030 25542
rect 13086 25540 13110 25542
rect 13166 25540 13190 25542
rect 13246 25540 13252 25542
rect 12944 25531 13252 25540
rect 13280 25498 13308 25706
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13188 24721 13216 24754
rect 13174 24712 13230 24721
rect 13174 24647 13230 24656
rect 12944 24508 13252 24517
rect 12944 24506 12950 24508
rect 13006 24506 13030 24508
rect 13086 24506 13110 24508
rect 13166 24506 13190 24508
rect 13246 24506 13252 24508
rect 13006 24454 13008 24506
rect 13188 24454 13190 24506
rect 12944 24452 12950 24454
rect 13006 24452 13030 24454
rect 13086 24452 13110 24454
rect 13166 24452 13190 24454
rect 13246 24452 13252 24454
rect 12944 24443 13252 24452
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 13188 23866 13216 24074
rect 13372 24070 13400 25978
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13280 23882 13308 24006
rect 13176 23860 13228 23866
rect 13280 23854 13400 23882
rect 13176 23802 13228 23808
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12716 23316 12768 23322
rect 12716 23258 12768 23264
rect 12624 23112 12676 23118
rect 12622 23080 12624 23089
rect 12676 23080 12678 23089
rect 12622 23015 12678 23024
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12636 22642 12664 22918
rect 12728 22642 12756 23258
rect 12820 22982 12848 23598
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 12944 23420 13252 23429
rect 12944 23418 12950 23420
rect 13006 23418 13030 23420
rect 13086 23418 13110 23420
rect 13166 23418 13190 23420
rect 13246 23418 13252 23420
rect 13006 23366 13008 23418
rect 13188 23366 13190 23418
rect 12944 23364 12950 23366
rect 13006 23364 13030 23366
rect 13086 23364 13110 23366
rect 13166 23364 13190 23366
rect 13246 23364 13252 23366
rect 12944 23355 13252 23364
rect 13280 23322 13308 23530
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 13004 22778 13032 22986
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12944 22332 13252 22341
rect 12944 22330 12950 22332
rect 13006 22330 13030 22332
rect 13086 22330 13110 22332
rect 13166 22330 13190 22332
rect 13246 22330 13252 22332
rect 13006 22278 13008 22330
rect 13188 22278 13190 22330
rect 12944 22276 12950 22278
rect 13006 22276 13030 22278
rect 13086 22276 13110 22278
rect 13166 22276 13190 22278
rect 13246 22276 13252 22278
rect 12944 22267 13252 22276
rect 12900 22228 12952 22234
rect 12254 21111 12310 21120
rect 12452 21134 12572 21162
rect 12728 22188 12900 22216
rect 12162 21040 12218 21049
rect 12162 20975 12218 20984
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12164 20868 12216 20874
rect 12164 20810 12216 20816
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12070 16960 12126 16969
rect 12070 16895 12126 16904
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11992 15366 12020 16186
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 12084 15094 12112 16895
rect 12072 15088 12124 15094
rect 11978 15056 12034 15065
rect 12072 15030 12124 15036
rect 11978 14991 11980 15000
rect 12032 14991 12034 15000
rect 11980 14962 12032 14968
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 11992 14793 12020 14826
rect 11978 14784 12034 14793
rect 11978 14719 12034 14728
rect 11978 14512 12034 14521
rect 11978 14447 11980 14456
rect 12032 14447 12034 14456
rect 11980 14418 12032 14424
rect 12084 14074 12112 14826
rect 12176 14618 12204 20810
rect 12268 20262 12296 20946
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12360 20369 12388 20402
rect 12346 20360 12402 20369
rect 12346 20295 12402 20304
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12268 19378 12296 20198
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12268 18834 12296 19110
rect 12360 18884 12388 19858
rect 12452 18952 12480 21134
rect 12532 20868 12584 20874
rect 12728 20856 12756 22188
rect 12900 22170 12952 22176
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12806 21584 12862 21593
rect 12806 21519 12862 21528
rect 12820 21026 12848 21519
rect 12912 21486 12940 21966
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13280 21486 13308 21830
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 12944 21244 13252 21253
rect 12944 21242 12950 21244
rect 13006 21242 13030 21244
rect 13086 21242 13110 21244
rect 13166 21242 13190 21244
rect 13246 21242 13252 21244
rect 13006 21190 13008 21242
rect 13188 21190 13190 21242
rect 12944 21188 12950 21190
rect 13006 21188 13030 21190
rect 13086 21188 13110 21190
rect 13166 21188 13190 21190
rect 13246 21188 13252 21190
rect 12944 21179 13252 21188
rect 12820 20998 12940 21026
rect 12912 20942 12940 20998
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12728 20828 12848 20856
rect 12532 20810 12584 20816
rect 12544 20505 12572 20810
rect 12530 20496 12586 20505
rect 12530 20431 12586 20440
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12636 20058 12664 20198
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 12544 19514 12572 19926
rect 12820 19922 12848 20828
rect 12944 20156 13252 20165
rect 12944 20154 12950 20156
rect 13006 20154 13030 20156
rect 13086 20154 13110 20156
rect 13166 20154 13190 20156
rect 13246 20154 13252 20156
rect 13006 20102 13008 20154
rect 13188 20102 13190 20154
rect 12944 20100 12950 20102
rect 13006 20100 13030 20102
rect 13086 20100 13110 20102
rect 13166 20100 13190 20102
rect 13246 20100 13252 20102
rect 12944 20091 13252 20100
rect 13082 19952 13138 19961
rect 12808 19916 12860 19922
rect 12860 19876 13032 19904
rect 13082 19887 13138 19896
rect 12808 19858 12860 19864
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 13004 19334 13032 19876
rect 13096 19378 13124 19887
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13280 19514 13308 19790
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 12728 19306 13032 19334
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13372 19334 13400 23854
rect 13464 22234 13492 27406
rect 13556 25838 13584 27814
rect 13636 27600 13688 27606
rect 13636 27542 13688 27548
rect 13648 25838 13676 27542
rect 13740 27062 13768 28698
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13832 28529 13860 28562
rect 13818 28520 13874 28529
rect 13818 28455 13874 28464
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13832 27441 13860 28086
rect 13924 27962 13952 30058
rect 14016 28762 14044 31726
rect 14096 31340 14148 31346
rect 14096 31282 14148 31288
rect 14004 28756 14056 28762
rect 14004 28698 14056 28704
rect 13924 27934 14044 27962
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13818 27432 13874 27441
rect 13818 27367 13874 27376
rect 13820 27328 13872 27334
rect 13820 27270 13872 27276
rect 13728 27056 13780 27062
rect 13728 26998 13780 27004
rect 13832 25906 13860 27270
rect 13924 26450 13952 27814
rect 14016 26874 14044 27934
rect 14108 27062 14136 31282
rect 14200 30410 14228 32302
rect 14292 32026 14320 32846
rect 14476 32348 14504 35006
rect 14556 35012 14608 35018
rect 14556 34954 14608 34960
rect 14568 33969 14596 34954
rect 14657 34844 14965 34853
rect 14657 34842 14663 34844
rect 14719 34842 14743 34844
rect 14799 34842 14823 34844
rect 14879 34842 14903 34844
rect 14959 34842 14965 34844
rect 14719 34790 14721 34842
rect 14901 34790 14903 34842
rect 14657 34788 14663 34790
rect 14719 34788 14743 34790
rect 14799 34788 14823 34790
rect 14879 34788 14903 34790
rect 14959 34788 14965 34790
rect 14657 34779 14965 34788
rect 14554 33960 14610 33969
rect 14554 33895 14610 33904
rect 14657 33756 14965 33765
rect 14657 33754 14663 33756
rect 14719 33754 14743 33756
rect 14799 33754 14823 33756
rect 14879 33754 14903 33756
rect 14959 33754 14965 33756
rect 14719 33702 14721 33754
rect 14901 33702 14903 33754
rect 14657 33700 14663 33702
rect 14719 33700 14743 33702
rect 14799 33700 14823 33702
rect 14879 33700 14903 33702
rect 14959 33700 14965 33702
rect 14657 33691 14965 33700
rect 14556 32836 14608 32842
rect 14556 32778 14608 32784
rect 14384 32320 14504 32348
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14292 30705 14320 31758
rect 14278 30696 14334 30705
rect 14278 30631 14334 30640
rect 14200 30382 14320 30410
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 14200 28540 14228 29106
rect 14292 28665 14320 30382
rect 14278 28656 14334 28665
rect 14278 28591 14334 28600
rect 14200 28512 14320 28540
rect 14188 27396 14240 27402
rect 14188 27338 14240 27344
rect 14096 27056 14148 27062
rect 14200 27033 14228 27338
rect 14096 26998 14148 27004
rect 14186 27024 14242 27033
rect 14186 26959 14242 26968
rect 14016 26846 14228 26874
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 14096 26784 14148 26790
rect 14096 26726 14148 26732
rect 13912 26444 13964 26450
rect 13912 26386 13964 26392
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13544 25832 13596 25838
rect 13636 25832 13688 25838
rect 13544 25774 13596 25780
rect 13634 25800 13636 25809
rect 13688 25800 13690 25809
rect 13556 25378 13584 25774
rect 13634 25735 13690 25744
rect 13556 25350 13676 25378
rect 13544 25220 13596 25226
rect 13544 25162 13596 25168
rect 13556 24410 13584 25162
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13556 23662 13584 24210
rect 13648 23662 13676 25350
rect 13912 25220 13964 25226
rect 13912 25162 13964 25168
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13556 22778 13584 23598
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13556 22545 13584 22578
rect 13542 22536 13598 22545
rect 13542 22471 13598 22480
rect 13648 22386 13676 23598
rect 13740 22574 13768 24006
rect 13832 23730 13860 24550
rect 13924 24177 13952 25162
rect 14016 24721 14044 26726
rect 14108 26042 14136 26726
rect 14096 26036 14148 26042
rect 14096 25978 14148 25984
rect 14200 25786 14228 26846
rect 14108 25758 14228 25786
rect 14002 24712 14058 24721
rect 14002 24647 14058 24656
rect 13910 24168 13966 24177
rect 13910 24103 13966 24112
rect 14108 24018 14136 25758
rect 14188 25696 14240 25702
rect 14186 25664 14188 25673
rect 14240 25664 14242 25673
rect 14186 25599 14242 25608
rect 14292 25514 14320 28512
rect 13924 23990 14136 24018
rect 14200 25486 14320 25514
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13820 22432 13872 22438
rect 13556 22358 13676 22386
rect 13726 22400 13782 22409
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 13464 19922 13492 21898
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13372 19306 13492 19334
rect 12452 18924 12618 18952
rect 12360 18856 12480 18884
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12268 14226 12296 18634
rect 12360 17610 12388 18702
rect 12452 18204 12480 18856
rect 12590 18816 12618 18924
rect 12590 18788 12664 18816
rect 12532 18216 12584 18222
rect 12452 18176 12532 18204
rect 12532 18158 12584 18164
rect 12438 18048 12494 18057
rect 12438 17983 12494 17992
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12452 16538 12480 17983
rect 12544 17377 12572 18158
rect 12530 17368 12586 17377
rect 12636 17338 12664 18788
rect 12728 18222 12756 19306
rect 12944 19068 13252 19077
rect 12944 19066 12950 19068
rect 13006 19066 13030 19068
rect 13086 19066 13110 19068
rect 13166 19066 13190 19068
rect 13246 19066 13252 19068
rect 13006 19014 13008 19066
rect 13188 19014 13190 19066
rect 12944 19012 12950 19014
rect 13006 19012 13030 19014
rect 13086 19012 13110 19014
rect 13166 19012 13190 19014
rect 13246 19012 13252 19014
rect 12944 19003 13252 19012
rect 12990 18864 13046 18873
rect 12990 18799 13046 18808
rect 13004 18766 13032 18799
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12530 17303 12586 17312
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12728 17218 12756 18158
rect 12636 17190 12756 17218
rect 12530 16824 12586 16833
rect 12530 16759 12532 16768
rect 12584 16759 12586 16768
rect 12532 16730 12584 16736
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12360 16510 12480 16538
rect 12360 16046 12388 16510
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16130 12480 16390
rect 12544 16250 12572 16594
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12636 16164 12664 17190
rect 12820 17066 12848 18158
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 12944 17980 13252 17989
rect 12944 17978 12950 17980
rect 13006 17978 13030 17980
rect 13086 17978 13110 17980
rect 13166 17978 13190 17980
rect 13246 17978 13252 17980
rect 13006 17926 13008 17978
rect 13188 17926 13190 17978
rect 12944 17924 12950 17926
rect 13006 17924 13030 17926
rect 13086 17924 13110 17926
rect 13166 17924 13190 17926
rect 13246 17924 13252 17926
rect 12944 17915 13252 17924
rect 13280 17882 13308 18090
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13372 17202 13400 18022
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 13188 17082 13216 17138
rect 13464 17134 13492 19306
rect 13556 18630 13584 22358
rect 13820 22374 13872 22380
rect 13726 22335 13782 22344
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 13648 21593 13676 22170
rect 13740 21690 13768 22335
rect 13832 22137 13860 22374
rect 13818 22128 13874 22137
rect 13818 22063 13874 22072
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13634 21584 13690 21593
rect 13924 21570 13952 23990
rect 14200 23882 14228 25486
rect 14384 24596 14412 32320
rect 14464 31952 14516 31958
rect 14464 31894 14516 31900
rect 14108 23854 14228 23882
rect 14292 24568 14412 24596
rect 14108 22094 14136 23854
rect 14188 23520 14240 23526
rect 14186 23488 14188 23497
rect 14240 23488 14242 23497
rect 14186 23423 14242 23432
rect 14292 23338 14320 24568
rect 13634 21519 13690 21528
rect 13740 21542 13952 21570
rect 14016 22066 14136 22094
rect 14200 23310 14320 23338
rect 13636 21480 13688 21486
rect 13636 21422 13688 21428
rect 13648 20806 13676 21422
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13648 18222 13676 19858
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13740 18170 13768 21542
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13832 21146 13860 21422
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13910 21040 13966 21049
rect 13832 20998 13910 21026
rect 13832 20058 13860 20998
rect 13910 20975 13966 20984
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13924 19961 13952 20538
rect 13910 19952 13966 19961
rect 13910 19887 13966 19896
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13832 19417 13860 19654
rect 13818 19408 13874 19417
rect 13818 19343 13874 19352
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13832 18766 13860 19246
rect 14016 18850 14044 22066
rect 14094 21584 14150 21593
rect 14094 21519 14150 21528
rect 14108 21078 14136 21519
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 14108 18873 14136 19110
rect 13924 18822 14044 18850
rect 14094 18864 14150 18873
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13820 18624 13872 18630
rect 13924 18601 13952 18822
rect 14094 18799 14150 18808
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13820 18566 13872 18572
rect 13910 18592 13966 18601
rect 13832 18290 13860 18566
rect 13910 18527 13966 18536
rect 13910 18320 13966 18329
rect 13820 18284 13872 18290
rect 13910 18255 13966 18264
rect 13820 18226 13872 18232
rect 13648 18034 13676 18158
rect 13740 18142 13860 18170
rect 13832 18086 13860 18142
rect 13820 18080 13872 18086
rect 13648 18006 13768 18034
rect 13820 18022 13872 18028
rect 13740 17762 13768 18006
rect 13818 17912 13874 17921
rect 13818 17847 13820 17856
rect 13872 17847 13874 17856
rect 13820 17818 13872 17824
rect 13544 17740 13596 17746
rect 13740 17734 13860 17762
rect 13544 17682 13596 17688
rect 13452 17128 13504 17134
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12716 16992 12768 16998
rect 12912 16980 12940 17070
rect 13188 17054 13308 17082
rect 13452 17070 13504 17076
rect 12878 16952 12940 16980
rect 12878 16946 12906 16952
rect 12716 16934 12768 16940
rect 12728 16266 12756 16934
rect 12820 16918 12906 16946
rect 12820 16590 12848 16918
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12944 16827 13252 16836
rect 12898 16688 12954 16697
rect 12898 16623 12954 16632
rect 12912 16590 12940 16623
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12900 16584 12952 16590
rect 13084 16584 13136 16590
rect 12900 16526 12952 16532
rect 13004 16544 13084 16572
rect 12820 16454 12848 16526
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 13004 16266 13032 16544
rect 13084 16526 13136 16532
rect 12728 16238 13032 16266
rect 12636 16136 12756 16164
rect 12452 16102 12572 16130
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12452 14890 12480 15914
rect 12544 14958 12572 16102
rect 12728 16096 12756 16136
rect 12636 16068 12756 16096
rect 12636 15162 12664 16068
rect 12808 16040 12860 16046
rect 12728 16000 12808 16028
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12728 14958 12756 16000
rect 12808 15982 12860 15988
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12532 14952 12584 14958
rect 12716 14952 12768 14958
rect 12532 14894 12584 14900
rect 12636 14912 12716 14940
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12636 14482 12664 14912
rect 12716 14894 12768 14900
rect 12714 14784 12770 14793
rect 12714 14719 12770 14728
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12176 14198 12296 14226
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12345 11836 12786
rect 11888 12436 11940 12442
rect 11992 12424 12020 13942
rect 12176 13138 12204 14198
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12268 13394 12296 14010
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12268 13297 12296 13330
rect 12254 13288 12310 13297
rect 12254 13223 12310 13232
rect 11940 12396 12020 12424
rect 11888 12378 11940 12384
rect 11794 12336 11850 12345
rect 11794 12271 11850 12280
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11256 10130 11284 10474
rect 11624 10130 11652 11018
rect 11716 10985 11744 11630
rect 11702 10976 11758 10985
rect 11702 10911 11758 10920
rect 11808 10742 11836 12038
rect 11886 11248 11942 11257
rect 11886 11183 11888 11192
rect 11940 11183 11942 11192
rect 11888 11154 11940 11160
rect 11992 11150 12020 12396
rect 12084 13110 12204 13138
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11980 10804 12032 10810
rect 11900 10764 11980 10792
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 11624 9654 11652 9862
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11520 9512 11572 9518
rect 11716 9500 11744 10406
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11572 9472 11744 9500
rect 11520 9454 11572 9460
rect 11256 9353 11284 9454
rect 11336 9376 11388 9382
rect 11242 9344 11298 9353
rect 11336 9318 11388 9324
rect 11242 9279 11298 9288
rect 11348 9178 11376 9318
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11440 9081 11468 9454
rect 11426 9072 11482 9081
rect 11426 9007 11482 9016
rect 11244 8968 11296 8974
rect 11150 8936 11206 8945
rect 11244 8910 11296 8916
rect 11150 8871 11206 8880
rect 11256 8820 11284 8910
rect 11164 8792 11284 8820
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10692 7404 10744 7410
rect 10796 7398 10916 7426
rect 10692 7346 10744 7352
rect 10888 7342 10916 7398
rect 11072 7342 11100 8230
rect 11164 7546 11192 8792
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 11624 8634 11652 9472
rect 11808 9353 11836 9998
rect 11900 9489 11928 10764
rect 11980 10746 12032 10752
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11886 9480 11942 9489
rect 11886 9415 11942 9424
rect 11794 9344 11850 9353
rect 11794 9279 11850 9288
rect 11702 9208 11758 9217
rect 11702 9143 11758 9152
rect 11716 8838 11744 9143
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11808 8634 11836 9046
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11518 8528 11574 8537
rect 11900 8498 11928 9415
rect 11992 9081 12020 9862
rect 11978 9072 12034 9081
rect 11978 9007 12034 9016
rect 11978 8936 12034 8945
rect 11978 8871 12034 8880
rect 11518 8463 11574 8472
rect 11888 8492 11940 8498
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11348 7857 11376 8298
rect 11440 7886 11468 8298
rect 11532 7954 11560 8463
rect 11888 8434 11940 8440
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11428 7880 11480 7886
rect 11334 7848 11390 7857
rect 11428 7822 11480 7828
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11334 7783 11390 7792
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10612 6304 10640 6802
rect 10692 6316 10744 6322
rect 10612 6276 10692 6304
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9784 5086 9904 5114
rect 9784 5030 9812 5086
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9876 4690 9904 5086
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 9968 2106 9996 5510
rect 10612 5370 10640 6276
rect 10692 6258 10744 6264
rect 10796 5778 10824 7142
rect 10888 6254 10916 7278
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10888 5642 10916 6190
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 11072 2774 11100 7278
rect 11624 7206 11652 7822
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6458 11192 6598
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 11808 4758 11836 7346
rect 11900 7002 11928 8026
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11992 5778 12020 8871
rect 12084 6866 12112 13110
rect 12254 12880 12310 12889
rect 12254 12815 12256 12824
rect 12308 12815 12310 12824
rect 12256 12786 12308 12792
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12176 11778 12204 12718
rect 12360 12238 12388 14350
rect 12530 13968 12586 13977
rect 12452 13926 12530 13954
rect 12452 12646 12480 13926
rect 12530 13903 12586 13912
rect 12636 13870 12664 14418
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13530 12572 13670
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12728 13410 12756 14719
rect 12820 13512 12848 15846
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 13280 15609 13308 17054
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13266 15600 13322 15609
rect 13266 15535 13322 15544
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13004 14929 13032 15438
rect 13096 15366 13124 15438
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13096 15201 13124 15302
rect 13082 15192 13138 15201
rect 13280 15162 13308 15438
rect 13082 15127 13138 15136
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 12990 14920 13046 14929
rect 12990 14855 13046 14864
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 12900 13524 12952 13530
rect 12820 13484 12900 13512
rect 12900 13466 12952 13472
rect 12728 13382 12848 13410
rect 12716 13320 12768 13326
rect 12622 13288 12678 13297
rect 12716 13262 12768 13268
rect 12622 13223 12678 13232
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12176 11750 12388 11778
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 10810 12204 11018
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12176 9625 12204 10542
rect 12268 10266 12296 11494
rect 12360 10792 12388 11750
rect 12360 10764 12480 10792
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12268 9761 12296 9862
rect 12254 9752 12310 9761
rect 12360 9704 12388 10610
rect 12452 10470 12480 10764
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12544 10282 12572 12718
rect 12636 11898 12664 13223
rect 12728 12442 12756 13262
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10606 12756 10950
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12254 9687 12310 9696
rect 12342 9676 12388 9704
rect 12452 10254 12572 10282
rect 12728 10266 12756 10542
rect 12624 10260 12676 10266
rect 12162 9616 12218 9625
rect 12218 9574 12296 9602
rect 12162 9551 12218 9560
rect 12268 7886 12296 9574
rect 12342 9466 12370 9676
rect 12452 9518 12480 10254
rect 12624 10202 12676 10208
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12636 9602 12664 10202
rect 12714 10160 12770 10169
rect 12820 10130 12848 13382
rect 13280 12714 13308 13670
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 13268 12232 13320 12238
rect 13266 12200 13268 12209
rect 13320 12200 13322 12209
rect 13266 12135 13322 12144
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 13280 11354 13308 11562
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12714 10095 12716 10104
rect 12768 10095 12770 10104
rect 12808 10124 12860 10130
rect 12716 10066 12768 10072
rect 12808 10066 12860 10072
rect 12806 10024 12862 10033
rect 12806 9959 12862 9968
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12544 9586 12664 9602
rect 12728 9586 12756 9862
rect 12532 9580 12664 9586
rect 12584 9574 12664 9580
rect 12716 9580 12768 9586
rect 12532 9522 12584 9528
rect 12716 9522 12768 9528
rect 12440 9512 12492 9518
rect 12342 9438 12388 9466
rect 12440 9454 12492 9460
rect 12360 9217 12388 9438
rect 12346 9208 12402 9217
rect 12346 9143 12402 9152
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8090 12388 8910
rect 12452 8566 12480 9454
rect 12714 8664 12770 8673
rect 12820 8650 12848 9959
rect 13004 9364 13032 10202
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12878 9336 13032 9364
rect 12878 9160 12906 9336
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 12878 9132 13032 9160
rect 12820 8622 12940 8650
rect 13004 8634 13032 9132
rect 12714 8599 12770 8608
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12624 8288 12676 8294
rect 12544 8248 12624 8276
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12256 7880 12308 7886
rect 12162 7848 12218 7857
rect 12256 7822 12308 7828
rect 12162 7783 12218 7792
rect 12176 7154 12204 7783
rect 12176 7126 12480 7154
rect 12346 6896 12402 6905
rect 12072 6860 12124 6866
rect 12346 6831 12402 6840
rect 12072 6802 12124 6808
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 5234 12020 5714
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 12176 4826 12204 6122
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 11808 4146 11836 4694
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 12360 3602 12388 6831
rect 12452 6474 12480 7126
rect 12544 6662 12572 8248
rect 12624 8230 12676 8236
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12452 6446 12572 6474
rect 12438 6352 12494 6361
rect 12544 6322 12572 6446
rect 12438 6287 12440 6296
rect 12492 6287 12494 6296
rect 12532 6316 12584 6322
rect 12440 6258 12492 6264
rect 12532 6258 12584 6264
rect 12636 5710 12664 7754
rect 12728 6848 12756 8599
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12820 8401 12848 8502
rect 12806 8392 12862 8401
rect 12806 8327 12862 8336
rect 12820 6984 12848 8327
rect 12912 8294 12940 8622
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 13280 7562 13308 9998
rect 13372 9602 13400 16934
rect 13556 16114 13584 17682
rect 13726 17504 13782 17513
rect 13726 17439 13782 17448
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13450 16008 13506 16017
rect 13450 15943 13506 15952
rect 13464 14618 13492 15943
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13648 14074 13676 17274
rect 13740 16522 13768 17439
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13726 16416 13782 16425
rect 13726 16351 13782 16360
rect 13740 14414 13768 16351
rect 13832 15586 13860 17734
rect 13924 17338 13952 18255
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14016 16946 14044 18702
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18426 14136 18566
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 14200 17513 14228 23310
rect 14370 23216 14426 23225
rect 14292 23174 14370 23202
rect 14292 22778 14320 23174
rect 14370 23151 14426 23160
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14278 22672 14334 22681
rect 14278 22607 14334 22616
rect 14292 22234 14320 22607
rect 14384 22438 14412 23054
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14476 22094 14504 31894
rect 14568 30841 14596 32778
rect 14657 32668 14965 32677
rect 14657 32666 14663 32668
rect 14719 32666 14743 32668
rect 14799 32666 14823 32668
rect 14879 32666 14903 32668
rect 14959 32666 14965 32668
rect 14719 32614 14721 32666
rect 14901 32614 14903 32666
rect 14657 32612 14663 32614
rect 14719 32612 14743 32614
rect 14799 32612 14823 32614
rect 14879 32612 14903 32614
rect 14959 32612 14965 32614
rect 14657 32603 14965 32612
rect 14657 31580 14965 31589
rect 14657 31578 14663 31580
rect 14719 31578 14743 31580
rect 14799 31578 14823 31580
rect 14879 31578 14903 31580
rect 14959 31578 14965 31580
rect 14719 31526 14721 31578
rect 14901 31526 14903 31578
rect 14657 31524 14663 31526
rect 14719 31524 14743 31526
rect 14799 31524 14823 31526
rect 14879 31524 14903 31526
rect 14959 31524 14965 31526
rect 14657 31515 14965 31524
rect 14554 30832 14610 30841
rect 14554 30767 14610 30776
rect 14657 30492 14965 30501
rect 14657 30490 14663 30492
rect 14719 30490 14743 30492
rect 14799 30490 14823 30492
rect 14879 30490 14903 30492
rect 14959 30490 14965 30492
rect 14719 30438 14721 30490
rect 14901 30438 14903 30490
rect 14657 30436 14663 30438
rect 14719 30436 14743 30438
rect 14799 30436 14823 30438
rect 14879 30436 14903 30438
rect 14959 30436 14965 30438
rect 14657 30427 14965 30436
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14568 25537 14596 29990
rect 14657 29404 14965 29413
rect 14657 29402 14663 29404
rect 14719 29402 14743 29404
rect 14799 29402 14823 29404
rect 14879 29402 14903 29404
rect 14959 29402 14965 29404
rect 14719 29350 14721 29402
rect 14901 29350 14903 29402
rect 14657 29348 14663 29350
rect 14719 29348 14743 29350
rect 14799 29348 14823 29350
rect 14879 29348 14903 29350
rect 14959 29348 14965 29350
rect 14657 29339 14965 29348
rect 14657 28316 14965 28325
rect 14657 28314 14663 28316
rect 14719 28314 14743 28316
rect 14799 28314 14823 28316
rect 14879 28314 14903 28316
rect 14959 28314 14965 28316
rect 14719 28262 14721 28314
rect 14901 28262 14903 28314
rect 14657 28260 14663 28262
rect 14719 28260 14743 28262
rect 14799 28260 14823 28262
rect 14879 28260 14903 28262
rect 14959 28260 14965 28262
rect 14657 28251 14965 28260
rect 14657 27228 14965 27237
rect 14657 27226 14663 27228
rect 14719 27226 14743 27228
rect 14799 27226 14823 27228
rect 14879 27226 14903 27228
rect 14959 27226 14965 27228
rect 14719 27174 14721 27226
rect 14901 27174 14903 27226
rect 14657 27172 14663 27174
rect 14719 27172 14743 27174
rect 14799 27172 14823 27174
rect 14879 27172 14903 27174
rect 14959 27172 14965 27174
rect 14657 27163 14965 27172
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14660 26761 14688 27066
rect 14646 26752 14702 26761
rect 14646 26687 14702 26696
rect 14657 26140 14965 26149
rect 14657 26138 14663 26140
rect 14719 26138 14743 26140
rect 14799 26138 14823 26140
rect 14879 26138 14903 26140
rect 14959 26138 14965 26140
rect 14719 26086 14721 26138
rect 14901 26086 14903 26138
rect 14657 26084 14663 26086
rect 14719 26084 14743 26086
rect 14799 26084 14823 26086
rect 14879 26084 14903 26086
rect 14959 26084 14965 26086
rect 14657 26075 14965 26084
rect 14554 25528 14610 25537
rect 14554 25463 14610 25472
rect 14556 25424 14608 25430
rect 14556 25366 14608 25372
rect 14384 22066 14504 22094
rect 14280 22024 14332 22030
rect 14384 22001 14412 22066
rect 14280 21966 14332 21972
rect 14370 21992 14426 22001
rect 14292 21434 14320 21966
rect 14370 21927 14426 21936
rect 14464 21480 14516 21486
rect 14292 21406 14412 21434
rect 14464 21422 14516 21428
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14292 21049 14320 21286
rect 14278 21040 14334 21049
rect 14278 20975 14334 20984
rect 14384 20346 14412 21406
rect 14292 20318 14412 20346
rect 14292 19334 14320 20318
rect 14370 20224 14426 20233
rect 14370 20159 14426 20168
rect 14384 19514 14412 20159
rect 14476 19514 14504 21422
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14464 19372 14516 19378
rect 14292 19306 14412 19334
rect 14464 19314 14516 19320
rect 14278 19136 14334 19145
rect 14278 19071 14334 19080
rect 14292 18970 14320 19071
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14186 17504 14242 17513
rect 14384 17490 14412 19306
rect 14476 18426 14504 19314
rect 14568 18766 14596 25366
rect 14657 25052 14965 25061
rect 14657 25050 14663 25052
rect 14719 25050 14743 25052
rect 14799 25050 14823 25052
rect 14879 25050 14903 25052
rect 14959 25050 14965 25052
rect 14719 24998 14721 25050
rect 14901 24998 14903 25050
rect 14657 24996 14663 24998
rect 14719 24996 14743 24998
rect 14799 24996 14823 24998
rect 14879 24996 14903 24998
rect 14959 24996 14965 24998
rect 14657 24987 14965 24996
rect 14657 23964 14965 23973
rect 14657 23962 14663 23964
rect 14719 23962 14743 23964
rect 14799 23962 14823 23964
rect 14879 23962 14903 23964
rect 14959 23962 14965 23964
rect 14719 23910 14721 23962
rect 14901 23910 14903 23962
rect 14657 23908 14663 23910
rect 14719 23908 14743 23910
rect 14799 23908 14823 23910
rect 14879 23908 14903 23910
rect 14959 23908 14965 23910
rect 14657 23899 14965 23908
rect 14657 22876 14965 22885
rect 14657 22874 14663 22876
rect 14719 22874 14743 22876
rect 14799 22874 14823 22876
rect 14879 22874 14903 22876
rect 14959 22874 14965 22876
rect 14719 22822 14721 22874
rect 14901 22822 14903 22874
rect 14657 22820 14663 22822
rect 14719 22820 14743 22822
rect 14799 22820 14823 22822
rect 14879 22820 14903 22822
rect 14959 22820 14965 22822
rect 14657 22811 14965 22820
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 14936 22506 14964 22714
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 14657 21788 14965 21797
rect 14657 21786 14663 21788
rect 14719 21786 14743 21788
rect 14799 21786 14823 21788
rect 14879 21786 14903 21788
rect 14959 21786 14965 21788
rect 14719 21734 14721 21786
rect 14901 21734 14903 21786
rect 14657 21732 14663 21734
rect 14719 21732 14743 21734
rect 14799 21732 14823 21734
rect 14879 21732 14903 21734
rect 14959 21732 14965 21734
rect 14657 21723 14965 21732
rect 14657 20700 14965 20709
rect 14657 20698 14663 20700
rect 14719 20698 14743 20700
rect 14799 20698 14823 20700
rect 14879 20698 14903 20700
rect 14959 20698 14965 20700
rect 14719 20646 14721 20698
rect 14901 20646 14903 20698
rect 14657 20644 14663 20646
rect 14719 20644 14743 20646
rect 14799 20644 14823 20646
rect 14879 20644 14903 20646
rect 14959 20644 14965 20646
rect 14657 20635 14965 20644
rect 14657 19612 14965 19621
rect 14657 19610 14663 19612
rect 14719 19610 14743 19612
rect 14799 19610 14823 19612
rect 14879 19610 14903 19612
rect 14959 19610 14965 19612
rect 14719 19558 14721 19610
rect 14901 19558 14903 19610
rect 14657 19556 14663 19558
rect 14719 19556 14743 19558
rect 14799 19556 14823 19558
rect 14879 19556 14903 19558
rect 14959 19556 14965 19558
rect 14657 19547 14965 19556
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14660 18612 14688 19450
rect 14568 18584 14688 18612
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14568 18034 14596 18584
rect 14657 18524 14965 18533
rect 14657 18522 14663 18524
rect 14719 18522 14743 18524
rect 14799 18522 14823 18524
rect 14879 18522 14903 18524
rect 14959 18522 14965 18524
rect 14719 18470 14721 18522
rect 14901 18470 14903 18522
rect 14657 18468 14663 18470
rect 14719 18468 14743 18470
rect 14799 18468 14823 18470
rect 14879 18468 14903 18470
rect 14959 18468 14965 18470
rect 14657 18459 14965 18468
rect 14186 17439 14242 17448
rect 14292 17462 14412 17490
rect 13924 16918 14044 16946
rect 13924 16726 13952 16918
rect 14292 16776 14320 17462
rect 14200 16748 14320 16776
rect 14372 16788 14424 16794
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 14200 16425 14228 16748
rect 14372 16730 14424 16736
rect 14278 16688 14334 16697
rect 14278 16623 14334 16632
rect 14292 16590 14320 16623
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14186 16416 14242 16425
rect 14186 16351 14242 16360
rect 14186 16144 14242 16153
rect 14186 16079 14242 16088
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15706 13952 15846
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13832 15558 14044 15586
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13726 13968 13782 13977
rect 13726 13903 13782 13912
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 13464 12442 13492 13398
rect 13740 13326 13768 13903
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13728 13184 13780 13190
rect 13648 13144 13728 13172
rect 13648 12968 13676 13144
rect 13728 13126 13780 13132
rect 13648 12940 13701 12968
rect 13673 12866 13701 12940
rect 13556 12850 13701 12866
rect 13832 12850 13860 14214
rect 14016 13802 14044 15558
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14108 15473 14136 15506
rect 14094 15464 14150 15473
rect 14094 15399 14150 15408
rect 14094 15328 14150 15337
rect 14094 15263 14150 15272
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 14108 13682 14136 15263
rect 14200 15094 14228 16079
rect 14384 15706 14412 16730
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14278 14784 14334 14793
rect 14278 14719 14334 14728
rect 14292 13938 14320 14719
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14186 13832 14242 13841
rect 14186 13767 14242 13776
rect 14280 13796 14332 13802
rect 14016 13654 14136 13682
rect 13910 12880 13966 12889
rect 13544 12844 13701 12850
rect 13596 12838 13701 12844
rect 13820 12844 13872 12850
rect 13544 12786 13596 12792
rect 13910 12815 13966 12824
rect 13820 12786 13872 12792
rect 13636 12776 13688 12782
rect 13688 12724 13701 12764
rect 13636 12718 13701 12724
rect 13673 12628 13701 12718
rect 13673 12600 13860 12628
rect 13924 12617 13952 12815
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13464 10130 13492 12174
rect 13832 12102 13860 12600
rect 13910 12608 13966 12617
rect 13910 12543 13966 12552
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13726 11928 13782 11937
rect 13636 11892 13688 11898
rect 13924 11898 13952 12378
rect 13726 11863 13782 11872
rect 13912 11892 13964 11898
rect 13636 11834 13688 11840
rect 13648 11762 13676 11834
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13634 10568 13690 10577
rect 13634 10503 13690 10512
rect 13648 10266 13676 10503
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13452 9716 13504 9722
rect 13504 9676 13676 9704
rect 13452 9658 13504 9664
rect 13372 9574 13584 9602
rect 13450 9480 13506 9489
rect 13450 9415 13506 9424
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13372 9178 13400 9318
rect 13464 9178 13492 9415
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13556 9110 13584 9574
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13556 8922 13584 9046
rect 13648 9042 13676 9676
rect 13740 9058 13768 11863
rect 13912 11834 13964 11840
rect 13910 11792 13966 11801
rect 13820 11756 13872 11762
rect 13910 11727 13966 11736
rect 13820 11698 13872 11704
rect 13832 10810 13860 11698
rect 13924 11354 13952 11727
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 14016 10266 14044 13654
rect 14200 13546 14228 13767
rect 14280 13738 14332 13744
rect 14108 13518 14228 13546
rect 14292 13530 14320 13738
rect 14384 13530 14412 14214
rect 14280 13524 14332 13530
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 13910 10160 13966 10169
rect 13910 10095 13966 10104
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 9353 13860 9454
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13636 9036 13688 9042
rect 13740 9030 13860 9058
rect 13636 8978 13688 8984
rect 13360 8900 13412 8906
rect 13556 8894 13676 8922
rect 13360 8842 13412 8848
rect 13372 7993 13400 8842
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 8294 13492 8774
rect 13464 8266 13584 8294
rect 13358 7984 13414 7993
rect 13358 7919 13414 7928
rect 13188 7546 13308 7562
rect 13176 7540 13308 7546
rect 13228 7534 13308 7540
rect 13176 7482 13228 7488
rect 13556 7478 13584 8266
rect 13648 7750 13676 8894
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7546 13676 7686
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13544 7472 13596 7478
rect 13740 7449 13768 8842
rect 13832 8378 13860 9030
rect 13924 8634 13952 10095
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13832 8350 13952 8378
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 8090 13860 8230
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13924 8022 13952 8350
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 14004 7472 14056 7478
rect 13544 7414 13596 7420
rect 13726 7440 13782 7449
rect 13452 7404 13504 7410
rect 14004 7414 14056 7420
rect 13726 7375 13782 7384
rect 13912 7404 13964 7410
rect 13452 7346 13504 7352
rect 13912 7346 13964 7352
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 13280 6984 13308 7278
rect 12820 6956 13032 6984
rect 12728 6820 12940 6848
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12728 6458 12756 6666
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12912 6361 12940 6820
rect 12898 6352 12954 6361
rect 12716 6316 12768 6322
rect 12898 6287 12954 6296
rect 12716 6258 12768 6264
rect 12728 5914 12756 6258
rect 13004 6236 13032 6956
rect 13096 6956 13308 6984
rect 13096 6440 13124 6956
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13096 6412 13308 6440
rect 12820 6208 13032 6236
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12820 5794 12848 6208
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 13280 5914 13308 6412
rect 13372 6390 13400 6666
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13372 5817 13400 6054
rect 12728 5766 12848 5794
rect 13358 5808 13414 5817
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12728 5234 12756 5766
rect 13358 5743 13414 5752
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12544 4622 12572 5170
rect 12820 4808 12848 5510
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 12820 4780 12940 4808
rect 12912 4622 12940 4780
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12544 4078 12572 4558
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12438 3496 12494 3505
rect 12438 3431 12494 3440
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 11072 2746 11192 2774
rect 11058 2680 11114 2689
rect 11058 2615 11114 2624
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 11072 2038 11100 2615
rect 8944 2032 8996 2038
rect 8944 1974 8996 1980
rect 11060 2032 11112 2038
rect 11060 1974 11112 1980
rect 7932 1964 7984 1970
rect 7932 1906 7984 1912
rect 8576 1964 8628 1970
rect 8576 1906 8628 1912
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 10140 1964 10192 1970
rect 10140 1906 10192 1912
rect 10876 1964 10928 1970
rect 10876 1906 10928 1912
rect 7380 1828 7432 1834
rect 7380 1770 7432 1776
rect 7944 1562 7972 1906
rect 8588 1562 8616 1906
rect 9324 1562 9352 1906
rect 9517 1660 9825 1669
rect 9517 1658 9523 1660
rect 9579 1658 9603 1660
rect 9659 1658 9683 1660
rect 9739 1658 9763 1660
rect 9819 1658 9825 1660
rect 9579 1606 9581 1658
rect 9761 1606 9763 1658
rect 9517 1604 9523 1606
rect 9579 1604 9603 1606
rect 9659 1604 9683 1606
rect 9739 1604 9763 1606
rect 9819 1604 9825 1606
rect 9517 1595 9825 1604
rect 10152 1562 10180 1906
rect 10888 1562 10916 1906
rect 11164 1902 11192 2746
rect 11794 2680 11850 2689
rect 11794 2615 11850 2624
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 11808 2106 11836 2615
rect 12452 2106 12480 3431
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 12440 2100 12492 2106
rect 12440 2042 12492 2048
rect 11612 1964 11664 1970
rect 11612 1906 11664 1912
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 11624 1562 11652 1906
rect 12360 1562 12388 1906
rect 5724 1556 5776 1562
rect 5724 1498 5776 1504
rect 6460 1556 6512 1562
rect 6460 1498 6512 1504
rect 7196 1556 7248 1562
rect 7196 1498 7248 1504
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 8576 1556 8628 1562
rect 8576 1498 8628 1504
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 10140 1556 10192 1562
rect 10140 1498 10192 1504
rect 10876 1556 10928 1562
rect 10876 1498 10928 1504
rect 11612 1556 11664 1562
rect 11612 1498 11664 1504
rect 12348 1556 12400 1562
rect 12348 1498 12400 1504
rect 12544 1426 12572 4014
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 13372 3670 13400 5646
rect 13464 4826 13492 7346
rect 13726 7168 13782 7177
rect 13726 7103 13782 7112
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13556 5370 13584 6802
rect 13634 6760 13690 6769
rect 13634 6695 13636 6704
rect 13688 6695 13690 6704
rect 13636 6666 13688 6672
rect 13740 5794 13768 7103
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13648 5766 13768 5794
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13648 3058 13676 5766
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13740 5273 13768 5578
rect 13726 5264 13782 5273
rect 13726 5199 13782 5208
rect 13832 3942 13860 6598
rect 13924 6254 13952 7346
rect 13912 6248 13964 6254
rect 13910 6216 13912 6225
rect 13964 6216 13966 6225
rect 13910 6151 13966 6160
rect 14016 5710 14044 7414
rect 14004 5704 14056 5710
rect 13910 5672 13966 5681
rect 14004 5646 14056 5652
rect 13910 5607 13966 5616
rect 13924 5574 13952 5607
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 14108 2774 14136 13518
rect 14280 13466 14332 13472
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14186 13424 14242 13433
rect 14476 13410 14504 18022
rect 14568 18006 14688 18034
rect 14554 17912 14610 17921
rect 14554 17847 14610 17856
rect 14568 17105 14596 17847
rect 14660 17746 14688 18006
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 14554 17096 14610 17105
rect 14554 17031 14610 17040
rect 14554 16960 14610 16969
rect 14554 16895 14610 16904
rect 14568 15502 14596 16895
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14186 13359 14242 13368
rect 14384 13382 14504 13410
rect 14200 12238 14228 13359
rect 14278 12880 14334 12889
rect 14278 12815 14334 12824
rect 14292 12374 14320 12815
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14278 12064 14334 12073
rect 14278 11999 14334 12008
rect 14186 11792 14242 11801
rect 14186 11727 14242 11736
rect 14200 11150 14228 11727
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14200 10441 14228 10610
rect 14186 10432 14242 10441
rect 14186 10367 14242 10376
rect 14292 10282 14320 11999
rect 14200 10254 14320 10282
rect 14200 7698 14228 10254
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9625 14320 9930
rect 14278 9616 14334 9625
rect 14278 9551 14334 9560
rect 14278 8256 14334 8265
rect 14278 8191 14334 8200
rect 14292 7886 14320 8191
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14200 7670 14320 7698
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14200 6089 14228 6394
rect 14186 6080 14242 6089
rect 14186 6015 14242 6024
rect 14292 5930 14320 7670
rect 14384 7546 14412 13382
rect 14462 12744 14518 12753
rect 14462 12679 14464 12688
rect 14516 12679 14518 12688
rect 14464 12650 14516 12656
rect 14568 12594 14596 14758
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 14646 13696 14702 13705
rect 14646 13631 14702 13640
rect 14660 13394 14688 13631
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 14476 12566 14596 12594
rect 14476 11354 14504 12566
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 14646 11520 14702 11529
rect 14646 11455 14702 11464
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14660 11218 14688 11455
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14738 6352 14794 6361
rect 14200 5902 14320 5930
rect 14200 5846 14228 5902
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14186 5672 14242 5681
rect 14186 5607 14242 5616
rect 14200 3534 14228 5607
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14384 3058 14412 6326
rect 14738 6287 14740 6296
rect 14792 6287 14794 6296
rect 14740 6258 14792 6264
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 15028 2774 15056 41386
rect 15108 37664 15160 37670
rect 15108 37606 15160 37612
rect 15120 37233 15148 37606
rect 15106 37224 15162 37233
rect 15106 37159 15162 37168
rect 15108 36032 15160 36038
rect 15106 36000 15108 36009
rect 15160 36000 15162 36009
rect 15106 35935 15162 35944
rect 15108 35556 15160 35562
rect 15108 35498 15160 35504
rect 15120 34921 15148 35498
rect 15106 34912 15162 34921
rect 15106 34847 15162 34856
rect 15108 32224 15160 32230
rect 15108 32166 15160 32172
rect 15120 30054 15148 32166
rect 15108 30048 15160 30054
rect 15108 29990 15160 29996
rect 15108 29028 15160 29034
rect 15108 28970 15160 28976
rect 15120 26217 15148 28970
rect 15106 26208 15162 26217
rect 15106 26143 15162 26152
rect 15108 24132 15160 24138
rect 15108 24074 15160 24080
rect 15120 24041 15148 24074
rect 15106 24032 15162 24041
rect 15106 23967 15162 23976
rect 15108 22976 15160 22982
rect 15106 22944 15108 22953
rect 15160 22944 15162 22953
rect 15106 22879 15162 22888
rect 15108 22840 15160 22846
rect 15108 22782 15160 22788
rect 15120 12434 15148 22782
rect 15212 22778 15240 42570
rect 15304 22914 15332 42638
rect 15384 37324 15436 37330
rect 15384 37266 15436 37272
rect 15396 35873 15424 37266
rect 15568 36100 15620 36106
rect 15568 36042 15620 36048
rect 15382 35864 15438 35873
rect 15382 35799 15438 35808
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 15382 34504 15438 34513
rect 15382 34439 15438 34448
rect 15396 33969 15424 34439
rect 15382 33960 15438 33969
rect 15382 33895 15438 33904
rect 15384 33516 15436 33522
rect 15384 33458 15436 33464
rect 15396 24596 15424 33458
rect 15488 31657 15516 35430
rect 15580 34513 15608 36042
rect 15660 34604 15712 34610
rect 15660 34546 15712 34552
rect 15566 34504 15622 34513
rect 15566 34439 15622 34448
rect 15568 32972 15620 32978
rect 15568 32914 15620 32920
rect 15580 32201 15608 32914
rect 15566 32192 15622 32201
rect 15566 32127 15622 32136
rect 15474 31648 15530 31657
rect 15474 31583 15530 31592
rect 15672 30569 15700 34546
rect 15752 31136 15804 31142
rect 15752 31078 15804 31084
rect 15658 30560 15714 30569
rect 15658 30495 15714 30504
rect 15568 30252 15620 30258
rect 15620 30212 15700 30240
rect 15568 30194 15620 30200
rect 15476 30184 15528 30190
rect 15476 30126 15528 30132
rect 15488 27577 15516 30126
rect 15568 30048 15620 30054
rect 15568 29990 15620 29996
rect 15580 28393 15608 29990
rect 15566 28384 15622 28393
rect 15566 28319 15622 28328
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15474 27568 15530 27577
rect 15474 27503 15530 27512
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15488 25945 15516 26182
rect 15474 25936 15530 25945
rect 15474 25871 15530 25880
rect 15580 25430 15608 28018
rect 15568 25424 15620 25430
rect 15568 25366 15620 25372
rect 15396 24568 15516 24596
rect 15292 22908 15344 22914
rect 15292 22850 15344 22856
rect 15488 22846 15516 24568
rect 15476 22840 15528 22846
rect 15476 22782 15528 22788
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15384 22704 15436 22710
rect 15672 22658 15700 30212
rect 15764 26246 15792 31078
rect 15844 27668 15896 27674
rect 15844 27610 15896 27616
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15856 23882 15884 27610
rect 15384 22646 15436 22652
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 15198 21856 15254 21865
rect 15198 21791 15254 21800
rect 15212 20602 15240 21791
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15212 17921 15240 19722
rect 15198 17912 15254 17921
rect 15198 17847 15254 17856
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 17513 15240 17614
rect 15198 17504 15254 17513
rect 15198 17439 15254 17448
rect 15200 17400 15252 17406
rect 15200 17342 15252 17348
rect 15212 14074 15240 17342
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15198 13152 15254 13161
rect 15198 13087 15254 13096
rect 15212 12986 15240 13087
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15120 12406 15240 12434
rect 15106 12064 15162 12073
rect 15106 11999 15162 12008
rect 15120 11150 15148 11999
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15106 10160 15162 10169
rect 15106 10095 15162 10104
rect 15120 8974 15148 10095
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15120 7721 15148 7754
rect 15106 7712 15162 7721
rect 15106 7647 15162 7656
rect 15212 6866 15240 12406
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15120 6633 15148 6666
rect 15106 6624 15162 6633
rect 15106 6559 15162 6568
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 5545 15148 5578
rect 15106 5536 15162 5545
rect 15106 5471 15162 5480
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 14108 2746 14228 2774
rect 15028 2746 15240 2774
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 14200 2106 14228 2746
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 14188 2100 14240 2106
rect 14188 2042 14240 2048
rect 13452 2032 13504 2038
rect 13452 1974 13504 1980
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 12944 1660 13252 1669
rect 12944 1658 12950 1660
rect 13006 1658 13030 1660
rect 13086 1658 13110 1660
rect 13166 1658 13190 1660
rect 13246 1658 13252 1660
rect 13006 1606 13008 1658
rect 13188 1606 13190 1658
rect 12944 1604 12950 1606
rect 13006 1604 13030 1606
rect 13086 1604 13110 1606
rect 13166 1604 13190 1606
rect 13246 1604 13252 1606
rect 12944 1595 13252 1604
rect 13280 1562 13308 1906
rect 13464 1562 13492 1974
rect 13728 1964 13780 1970
rect 13728 1906 13780 1912
rect 13740 1562 13768 1906
rect 15212 1902 15240 2746
rect 15200 1896 15252 1902
rect 15200 1838 15252 1844
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 13452 1556 13504 1562
rect 13452 1498 13504 1504
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 12532 1420 12584 1426
rect 12532 1362 12584 1368
rect 15304 1358 15332 22442
rect 15396 1902 15424 22646
rect 15488 22630 15700 22658
rect 15764 23854 15884 23882
rect 15488 19786 15516 22630
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15474 19680 15530 19689
rect 15474 19615 15530 19624
rect 15488 17338 15516 19615
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15488 14521 15516 16050
rect 15474 14512 15530 14521
rect 15474 14447 15530 14456
rect 15474 14104 15530 14113
rect 15474 14039 15530 14048
rect 15488 12238 15516 14039
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15580 11898 15608 22374
rect 15672 15994 15700 22510
rect 15764 16114 15792 23854
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15672 15966 15792 15994
rect 15658 15872 15714 15881
rect 15658 15807 15714 15816
rect 15672 13326 15700 15807
rect 15764 15502 15792 15966
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15856 13190 15884 21898
rect 15948 21486 15976 22578
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15936 20732 15988 20738
rect 15936 20674 15988 20680
rect 15948 17406 15976 20674
rect 15936 17400 15988 17406
rect 15936 17342 15988 17348
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15856 10946 15884 13126
rect 15948 12442 15976 16050
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15844 10940 15896 10946
rect 15844 10882 15896 10888
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 9897 15516 10406
rect 15474 9888 15530 9897
rect 15474 9823 15530 9832
rect 15384 1896 15436 1902
rect 15384 1838 15436 1844
rect 3792 1352 3844 1358
rect 4620 1352 4672 1358
rect 3792 1294 3844 1300
rect 4618 1320 4620 1329
rect 5356 1352 5408 1358
rect 4672 1320 4674 1329
rect 2778 54 3096 82
rect 3514 82 3570 160
rect 3804 82 3832 1294
rect 4252 1284 4304 1290
rect 5354 1320 5356 1329
rect 5724 1352 5776 1358
rect 5408 1320 5410 1329
rect 4618 1255 4674 1264
rect 5172 1284 5224 1290
rect 4252 1226 4304 1232
rect 5724 1294 5776 1300
rect 6460 1352 6512 1358
rect 6460 1294 6512 1300
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 10140 1352 10192 1358
rect 10140 1294 10192 1300
rect 10876 1352 10928 1358
rect 10876 1294 10928 1300
rect 11612 1352 11664 1358
rect 11612 1294 11664 1300
rect 12348 1352 12400 1358
rect 12348 1294 12400 1300
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 13912 1352 13964 1358
rect 13912 1294 13964 1300
rect 14556 1352 14608 1358
rect 14556 1294 14608 1300
rect 15292 1352 15344 1358
rect 15292 1294 15344 1300
rect 5354 1255 5410 1264
rect 5172 1226 5224 1232
rect 4264 160 4292 1226
rect 4376 1116 4684 1125
rect 4376 1114 4382 1116
rect 4438 1114 4462 1116
rect 4518 1114 4542 1116
rect 4598 1114 4622 1116
rect 4678 1114 4684 1116
rect 4438 1062 4440 1114
rect 4620 1062 4622 1114
rect 4376 1060 4382 1062
rect 4438 1060 4462 1062
rect 4518 1060 4542 1062
rect 4598 1060 4622 1062
rect 4678 1060 4684 1062
rect 4376 1051 4684 1060
rect 3514 54 3832 82
rect 2778 0 2834 54
rect 3514 0 3570 54
rect 4250 0 4306 160
rect 4986 82 5042 160
rect 5184 82 5212 1226
rect 5736 160 5764 1294
rect 6472 160 6500 1294
rect 7208 160 7236 1294
rect 7803 1116 8111 1125
rect 7803 1114 7809 1116
rect 7865 1114 7889 1116
rect 7945 1114 7969 1116
rect 8025 1114 8049 1116
rect 8105 1114 8111 1116
rect 7865 1062 7867 1114
rect 8047 1062 8049 1114
rect 7803 1060 7809 1062
rect 7865 1060 7889 1062
rect 7945 1060 7969 1062
rect 8025 1060 8049 1062
rect 8105 1060 8111 1062
rect 7803 1051 8111 1060
rect 7944 190 8064 218
rect 7944 160 7972 190
rect 4986 54 5212 82
rect 4986 0 5042 54
rect 5722 0 5778 160
rect 6458 0 6514 160
rect 7194 0 7250 160
rect 7930 0 7986 160
rect 8036 82 8064 190
rect 8220 82 8248 1294
rect 8680 160 8708 1294
rect 8036 54 8248 82
rect 8666 0 8722 160
rect 9402 82 9458 160
rect 9692 82 9720 1294
rect 10152 160 10180 1294
rect 10888 160 10916 1294
rect 11230 1116 11538 1125
rect 11230 1114 11236 1116
rect 11292 1114 11316 1116
rect 11372 1114 11396 1116
rect 11452 1114 11476 1116
rect 11532 1114 11538 1116
rect 11292 1062 11294 1114
rect 11474 1062 11476 1114
rect 11230 1060 11236 1062
rect 11292 1060 11316 1062
rect 11372 1060 11396 1062
rect 11452 1060 11476 1062
rect 11532 1060 11538 1062
rect 11230 1051 11538 1060
rect 11624 160 11652 1294
rect 12360 160 12388 1294
rect 13096 190 13216 218
rect 13096 160 13124 190
rect 9402 54 9720 82
rect 9402 0 9458 54
rect 10138 0 10194 160
rect 10874 0 10930 160
rect 11610 0 11666 160
rect 12346 0 12402 160
rect 13082 0 13138 160
rect 13188 82 13216 190
rect 13372 82 13400 1294
rect 13188 54 13400 82
rect 13818 82 13874 160
rect 13924 82 13952 1294
rect 14568 160 14596 1294
rect 15292 1216 15344 1222
rect 15292 1158 15344 1164
rect 14657 1116 14965 1125
rect 14657 1114 14663 1116
rect 14719 1114 14743 1116
rect 14799 1114 14823 1116
rect 14879 1114 14903 1116
rect 14959 1114 14965 1116
rect 14719 1062 14721 1114
rect 14901 1062 14903 1114
rect 14657 1060 14663 1062
rect 14719 1060 14743 1062
rect 14799 1060 14823 1062
rect 14879 1060 14903 1062
rect 14959 1060 14965 1062
rect 14657 1051 14965 1060
rect 15304 160 15332 1158
rect 13818 54 13952 82
rect 13818 0 13874 54
rect 14554 0 14610 160
rect 15290 0 15346 160
<< via2 >>
rect 4382 43546 4438 43548
rect 4462 43546 4518 43548
rect 4542 43546 4598 43548
rect 4622 43546 4678 43548
rect 4382 43494 4428 43546
rect 4428 43494 4438 43546
rect 4462 43494 4492 43546
rect 4492 43494 4504 43546
rect 4504 43494 4518 43546
rect 4542 43494 4556 43546
rect 4556 43494 4568 43546
rect 4568 43494 4598 43546
rect 4622 43494 4632 43546
rect 4632 43494 4678 43546
rect 4382 43492 4438 43494
rect 4462 43492 4518 43494
rect 4542 43492 4598 43494
rect 4622 43492 4678 43494
rect 7809 43546 7865 43548
rect 7889 43546 7945 43548
rect 7969 43546 8025 43548
rect 8049 43546 8105 43548
rect 7809 43494 7855 43546
rect 7855 43494 7865 43546
rect 7889 43494 7919 43546
rect 7919 43494 7931 43546
rect 7931 43494 7945 43546
rect 7969 43494 7983 43546
rect 7983 43494 7995 43546
rect 7995 43494 8025 43546
rect 8049 43494 8059 43546
rect 8059 43494 8105 43546
rect 7809 43492 7865 43494
rect 7889 43492 7945 43494
rect 7969 43492 8025 43494
rect 8049 43492 8105 43494
rect 11236 43546 11292 43548
rect 11316 43546 11372 43548
rect 11396 43546 11452 43548
rect 11476 43546 11532 43548
rect 11236 43494 11282 43546
rect 11282 43494 11292 43546
rect 11316 43494 11346 43546
rect 11346 43494 11358 43546
rect 11358 43494 11372 43546
rect 11396 43494 11410 43546
rect 11410 43494 11422 43546
rect 11422 43494 11452 43546
rect 11476 43494 11486 43546
rect 11486 43494 11532 43546
rect 11236 43492 11292 43494
rect 11316 43492 11372 43494
rect 11396 43492 11452 43494
rect 11476 43492 11532 43494
rect 754 40840 810 40896
rect 754 40024 810 40080
rect 754 39208 810 39264
rect 754 37576 810 37632
rect 754 36760 810 36816
rect 754 35944 810 36000
rect 754 35128 810 35184
rect 754 33496 810 33552
rect 754 32680 810 32736
rect 754 31864 810 31920
rect 754 31048 810 31104
rect 754 29416 810 29472
rect 754 27784 810 27840
rect 754 26968 810 27024
rect 754 25336 810 25392
rect 754 24520 810 24576
rect 754 23704 810 23760
rect 754 22888 810 22944
rect 754 22072 810 22128
rect 754 21256 810 21312
rect 754 19624 810 19680
rect 754 17992 810 18048
rect 754 17176 810 17232
rect 754 15544 810 15600
rect 846 14764 848 14784
rect 848 14764 900 14784
rect 900 14764 902 14784
rect 846 14728 902 14764
rect 846 13912 902 13968
rect 846 13132 848 13152
rect 848 13132 900 13152
rect 900 13132 902 13152
rect 846 13096 902 13132
rect 846 12280 902 12336
rect 1398 38528 1454 38584
rect 2669 43002 2725 43004
rect 2749 43002 2805 43004
rect 2829 43002 2885 43004
rect 2909 43002 2965 43004
rect 2669 42950 2715 43002
rect 2715 42950 2725 43002
rect 2749 42950 2779 43002
rect 2779 42950 2791 43002
rect 2791 42950 2805 43002
rect 2829 42950 2843 43002
rect 2843 42950 2855 43002
rect 2855 42950 2885 43002
rect 2909 42950 2919 43002
rect 2919 42950 2965 43002
rect 2669 42948 2725 42950
rect 2749 42948 2805 42950
rect 2829 42948 2885 42950
rect 2909 42948 2965 42950
rect 1398 34448 1454 34504
rect 2669 41914 2725 41916
rect 2749 41914 2805 41916
rect 2829 41914 2885 41916
rect 2909 41914 2965 41916
rect 2669 41862 2715 41914
rect 2715 41862 2725 41914
rect 2749 41862 2779 41914
rect 2779 41862 2791 41914
rect 2791 41862 2805 41914
rect 2829 41862 2843 41914
rect 2843 41862 2855 41914
rect 2855 41862 2885 41914
rect 2909 41862 2919 41914
rect 2919 41862 2965 41914
rect 2669 41860 2725 41862
rect 2749 41860 2805 41862
rect 2829 41860 2885 41862
rect 2909 41860 2965 41862
rect 2669 40826 2725 40828
rect 2749 40826 2805 40828
rect 2829 40826 2885 40828
rect 2909 40826 2965 40828
rect 2669 40774 2715 40826
rect 2715 40774 2725 40826
rect 2749 40774 2779 40826
rect 2779 40774 2791 40826
rect 2791 40774 2805 40826
rect 2829 40774 2843 40826
rect 2843 40774 2855 40826
rect 2855 40774 2885 40826
rect 2909 40774 2919 40826
rect 2919 40774 2965 40826
rect 2669 40772 2725 40774
rect 2749 40772 2805 40774
rect 2829 40772 2885 40774
rect 2909 40772 2965 40774
rect 2669 39738 2725 39740
rect 2749 39738 2805 39740
rect 2829 39738 2885 39740
rect 2909 39738 2965 39740
rect 2669 39686 2715 39738
rect 2715 39686 2725 39738
rect 2749 39686 2779 39738
rect 2779 39686 2791 39738
rect 2791 39686 2805 39738
rect 2829 39686 2843 39738
rect 2843 39686 2855 39738
rect 2855 39686 2885 39738
rect 2909 39686 2919 39738
rect 2919 39686 2965 39738
rect 2669 39684 2725 39686
rect 2749 39684 2805 39686
rect 2829 39684 2885 39686
rect 2909 39684 2965 39686
rect 2669 38650 2725 38652
rect 2749 38650 2805 38652
rect 2829 38650 2885 38652
rect 2909 38650 2965 38652
rect 2669 38598 2715 38650
rect 2715 38598 2725 38650
rect 2749 38598 2779 38650
rect 2779 38598 2791 38650
rect 2791 38598 2805 38650
rect 2829 38598 2843 38650
rect 2843 38598 2855 38650
rect 2855 38598 2885 38650
rect 2909 38598 2919 38650
rect 2919 38598 2965 38650
rect 2669 38596 2725 38598
rect 2749 38596 2805 38598
rect 2829 38596 2885 38598
rect 2909 38596 2965 38598
rect 2669 37562 2725 37564
rect 2749 37562 2805 37564
rect 2829 37562 2885 37564
rect 2909 37562 2965 37564
rect 2669 37510 2715 37562
rect 2715 37510 2725 37562
rect 2749 37510 2779 37562
rect 2779 37510 2791 37562
rect 2791 37510 2805 37562
rect 2829 37510 2843 37562
rect 2843 37510 2855 37562
rect 2855 37510 2885 37562
rect 2909 37510 2919 37562
rect 2919 37510 2965 37562
rect 2669 37508 2725 37510
rect 2749 37508 2805 37510
rect 2829 37508 2885 37510
rect 2909 37508 2965 37510
rect 2669 36474 2725 36476
rect 2749 36474 2805 36476
rect 2829 36474 2885 36476
rect 2909 36474 2965 36476
rect 2669 36422 2715 36474
rect 2715 36422 2725 36474
rect 2749 36422 2779 36474
rect 2779 36422 2791 36474
rect 2791 36422 2805 36474
rect 2829 36422 2843 36474
rect 2843 36422 2855 36474
rect 2855 36422 2885 36474
rect 2909 36422 2919 36474
rect 2919 36422 2965 36474
rect 2669 36420 2725 36422
rect 2749 36420 2805 36422
rect 2829 36420 2885 36422
rect 2909 36420 2965 36422
rect 2669 35386 2725 35388
rect 2749 35386 2805 35388
rect 2829 35386 2885 35388
rect 2909 35386 2965 35388
rect 2669 35334 2715 35386
rect 2715 35334 2725 35386
rect 2749 35334 2779 35386
rect 2779 35334 2791 35386
rect 2791 35334 2805 35386
rect 2829 35334 2843 35386
rect 2843 35334 2855 35386
rect 2855 35334 2885 35386
rect 2909 35334 2919 35386
rect 2919 35334 2965 35386
rect 2669 35332 2725 35334
rect 2749 35332 2805 35334
rect 2829 35332 2885 35334
rect 2909 35332 2965 35334
rect 2669 34298 2725 34300
rect 2749 34298 2805 34300
rect 2829 34298 2885 34300
rect 2909 34298 2965 34300
rect 2669 34246 2715 34298
rect 2715 34246 2725 34298
rect 2749 34246 2779 34298
rect 2779 34246 2791 34298
rect 2791 34246 2805 34298
rect 2829 34246 2843 34298
rect 2843 34246 2855 34298
rect 2855 34246 2885 34298
rect 2909 34246 2919 34298
rect 2919 34246 2965 34298
rect 2669 34244 2725 34246
rect 2749 34244 2805 34246
rect 2829 34244 2885 34246
rect 2909 34244 2965 34246
rect 2669 33210 2725 33212
rect 2749 33210 2805 33212
rect 2829 33210 2885 33212
rect 2909 33210 2965 33212
rect 2669 33158 2715 33210
rect 2715 33158 2725 33210
rect 2749 33158 2779 33210
rect 2779 33158 2791 33210
rect 2791 33158 2805 33210
rect 2829 33158 2843 33210
rect 2843 33158 2855 33210
rect 2855 33158 2885 33210
rect 2909 33158 2919 33210
rect 2919 33158 2965 33210
rect 2669 33156 2725 33158
rect 2749 33156 2805 33158
rect 2829 33156 2885 33158
rect 2909 33156 2965 33158
rect 1398 30232 1454 30288
rect 1398 28872 1454 28928
rect 846 11500 848 11520
rect 848 11500 900 11520
rect 900 11500 902 11520
rect 846 11464 902 11500
rect 1030 9832 1086 9888
rect 1490 26152 1546 26208
rect 1398 20576 1454 20632
rect 1490 19216 1546 19272
rect 1490 16496 1546 16552
rect 1674 23160 1730 23216
rect 1674 19216 1730 19272
rect 1582 10956 1584 10976
rect 1584 10956 1636 10976
rect 1636 10956 1638 10976
rect 1582 10920 1638 10956
rect 1582 9560 1638 9616
rect 1766 9580 1822 9616
rect 1766 9560 1768 9580
rect 1768 9560 1820 9580
rect 1820 9560 1822 9580
rect 2669 32122 2725 32124
rect 2749 32122 2805 32124
rect 2829 32122 2885 32124
rect 2909 32122 2965 32124
rect 2669 32070 2715 32122
rect 2715 32070 2725 32122
rect 2749 32070 2779 32122
rect 2779 32070 2791 32122
rect 2791 32070 2805 32122
rect 2829 32070 2843 32122
rect 2843 32070 2855 32122
rect 2855 32070 2885 32122
rect 2909 32070 2919 32122
rect 2919 32070 2965 32122
rect 2669 32068 2725 32070
rect 2749 32068 2805 32070
rect 2829 32068 2885 32070
rect 2909 32068 2965 32070
rect 2669 31034 2725 31036
rect 2749 31034 2805 31036
rect 2829 31034 2885 31036
rect 2909 31034 2965 31036
rect 2669 30982 2715 31034
rect 2715 30982 2725 31034
rect 2749 30982 2779 31034
rect 2779 30982 2791 31034
rect 2791 30982 2805 31034
rect 2829 30982 2843 31034
rect 2843 30982 2855 31034
rect 2855 30982 2885 31034
rect 2909 30982 2919 31034
rect 2919 30982 2965 31034
rect 2669 30980 2725 30982
rect 2749 30980 2805 30982
rect 2829 30980 2885 30982
rect 2909 30980 2965 30982
rect 2669 29946 2725 29948
rect 2749 29946 2805 29948
rect 2829 29946 2885 29948
rect 2909 29946 2965 29948
rect 2669 29894 2715 29946
rect 2715 29894 2725 29946
rect 2749 29894 2779 29946
rect 2779 29894 2791 29946
rect 2791 29894 2805 29946
rect 2829 29894 2843 29946
rect 2843 29894 2855 29946
rect 2855 29894 2885 29946
rect 2909 29894 2919 29946
rect 2919 29894 2965 29946
rect 2669 29892 2725 29894
rect 2749 29892 2805 29894
rect 2829 29892 2885 29894
rect 2909 29892 2965 29894
rect 1950 20304 2006 20360
rect 2669 28858 2725 28860
rect 2749 28858 2805 28860
rect 2829 28858 2885 28860
rect 2909 28858 2965 28860
rect 2669 28806 2715 28858
rect 2715 28806 2725 28858
rect 2749 28806 2779 28858
rect 2779 28806 2791 28858
rect 2791 28806 2805 28858
rect 2829 28806 2843 28858
rect 2843 28806 2855 28858
rect 2855 28806 2885 28858
rect 2909 28806 2919 28858
rect 2919 28806 2965 28858
rect 2669 28804 2725 28806
rect 2749 28804 2805 28806
rect 2829 28804 2885 28806
rect 2909 28804 2965 28806
rect 2669 27770 2725 27772
rect 2749 27770 2805 27772
rect 2829 27770 2885 27772
rect 2909 27770 2965 27772
rect 2669 27718 2715 27770
rect 2715 27718 2725 27770
rect 2749 27718 2779 27770
rect 2779 27718 2791 27770
rect 2791 27718 2805 27770
rect 2829 27718 2843 27770
rect 2843 27718 2855 27770
rect 2855 27718 2885 27770
rect 2909 27718 2919 27770
rect 2919 27718 2965 27770
rect 2669 27716 2725 27718
rect 2749 27716 2805 27718
rect 2829 27716 2885 27718
rect 2909 27716 2965 27718
rect 6096 43002 6152 43004
rect 6176 43002 6232 43004
rect 6256 43002 6312 43004
rect 6336 43002 6392 43004
rect 6096 42950 6142 43002
rect 6142 42950 6152 43002
rect 6176 42950 6206 43002
rect 6206 42950 6218 43002
rect 6218 42950 6232 43002
rect 6256 42950 6270 43002
rect 6270 42950 6282 43002
rect 6282 42950 6312 43002
rect 6336 42950 6346 43002
rect 6346 42950 6392 43002
rect 6096 42948 6152 42950
rect 6176 42948 6232 42950
rect 6256 42948 6312 42950
rect 6336 42948 6392 42950
rect 9523 43002 9579 43004
rect 9603 43002 9659 43004
rect 9683 43002 9739 43004
rect 9763 43002 9819 43004
rect 9523 42950 9569 43002
rect 9569 42950 9579 43002
rect 9603 42950 9633 43002
rect 9633 42950 9645 43002
rect 9645 42950 9659 43002
rect 9683 42950 9697 43002
rect 9697 42950 9709 43002
rect 9709 42950 9739 43002
rect 9763 42950 9773 43002
rect 9773 42950 9819 43002
rect 9523 42948 9579 42950
rect 9603 42948 9659 42950
rect 9683 42948 9739 42950
rect 9763 42948 9819 42950
rect 12950 43002 13006 43004
rect 13030 43002 13086 43004
rect 13110 43002 13166 43004
rect 13190 43002 13246 43004
rect 12950 42950 12996 43002
rect 12996 42950 13006 43002
rect 13030 42950 13060 43002
rect 13060 42950 13072 43002
rect 13072 42950 13086 43002
rect 13110 42950 13124 43002
rect 13124 42950 13136 43002
rect 13136 42950 13166 43002
rect 13190 42950 13200 43002
rect 13200 42950 13246 43002
rect 12950 42948 13006 42950
rect 13030 42948 13086 42950
rect 13110 42948 13166 42950
rect 13190 42948 13246 42950
rect 2669 26682 2725 26684
rect 2749 26682 2805 26684
rect 2829 26682 2885 26684
rect 2909 26682 2965 26684
rect 2669 26630 2715 26682
rect 2715 26630 2725 26682
rect 2749 26630 2779 26682
rect 2779 26630 2791 26682
rect 2791 26630 2805 26682
rect 2829 26630 2843 26682
rect 2843 26630 2855 26682
rect 2855 26630 2885 26682
rect 2909 26630 2919 26682
rect 2919 26630 2965 26682
rect 2669 26628 2725 26630
rect 2749 26628 2805 26630
rect 2829 26628 2885 26630
rect 2909 26628 2965 26630
rect 2669 25594 2725 25596
rect 2749 25594 2805 25596
rect 2829 25594 2885 25596
rect 2909 25594 2965 25596
rect 2669 25542 2715 25594
rect 2715 25542 2725 25594
rect 2749 25542 2779 25594
rect 2779 25542 2791 25594
rect 2791 25542 2805 25594
rect 2829 25542 2843 25594
rect 2843 25542 2855 25594
rect 2855 25542 2885 25594
rect 2909 25542 2919 25594
rect 2919 25542 2965 25594
rect 2669 25540 2725 25542
rect 2749 25540 2805 25542
rect 2829 25540 2885 25542
rect 2909 25540 2965 25542
rect 2669 24506 2725 24508
rect 2749 24506 2805 24508
rect 2829 24506 2885 24508
rect 2909 24506 2965 24508
rect 2669 24454 2715 24506
rect 2715 24454 2725 24506
rect 2749 24454 2779 24506
rect 2779 24454 2791 24506
rect 2791 24454 2805 24506
rect 2829 24454 2843 24506
rect 2843 24454 2855 24506
rect 2855 24454 2885 24506
rect 2909 24454 2919 24506
rect 2919 24454 2965 24506
rect 2669 24452 2725 24454
rect 2749 24452 2805 24454
rect 2829 24452 2885 24454
rect 2909 24452 2965 24454
rect 2669 23418 2725 23420
rect 2749 23418 2805 23420
rect 2829 23418 2885 23420
rect 2909 23418 2965 23420
rect 2669 23366 2715 23418
rect 2715 23366 2725 23418
rect 2749 23366 2779 23418
rect 2779 23366 2791 23418
rect 2791 23366 2805 23418
rect 2829 23366 2843 23418
rect 2843 23366 2855 23418
rect 2855 23366 2885 23418
rect 2909 23366 2919 23418
rect 2919 23366 2965 23418
rect 2669 23364 2725 23366
rect 2749 23364 2805 23366
rect 2829 23364 2885 23366
rect 2909 23364 2965 23366
rect 2669 22330 2725 22332
rect 2749 22330 2805 22332
rect 2829 22330 2885 22332
rect 2909 22330 2965 22332
rect 2669 22278 2715 22330
rect 2715 22278 2725 22330
rect 2749 22278 2779 22330
rect 2779 22278 2791 22330
rect 2791 22278 2805 22330
rect 2829 22278 2843 22330
rect 2843 22278 2855 22330
rect 2855 22278 2885 22330
rect 2909 22278 2919 22330
rect 2919 22278 2965 22330
rect 2669 22276 2725 22278
rect 2749 22276 2805 22278
rect 2829 22276 2885 22278
rect 2909 22276 2965 22278
rect 2669 21242 2725 21244
rect 2749 21242 2805 21244
rect 2829 21242 2885 21244
rect 2909 21242 2965 21244
rect 2669 21190 2715 21242
rect 2715 21190 2725 21242
rect 2749 21190 2779 21242
rect 2779 21190 2791 21242
rect 2791 21190 2805 21242
rect 2829 21190 2843 21242
rect 2843 21190 2855 21242
rect 2855 21190 2885 21242
rect 2909 21190 2919 21242
rect 2919 21190 2965 21242
rect 2669 21188 2725 21190
rect 2749 21188 2805 21190
rect 2829 21188 2885 21190
rect 2909 21188 2965 21190
rect 2669 20154 2725 20156
rect 2749 20154 2805 20156
rect 2829 20154 2885 20156
rect 2909 20154 2965 20156
rect 2669 20102 2715 20154
rect 2715 20102 2725 20154
rect 2749 20102 2779 20154
rect 2779 20102 2791 20154
rect 2791 20102 2805 20154
rect 2829 20102 2843 20154
rect 2843 20102 2855 20154
rect 2855 20102 2885 20154
rect 2909 20102 2919 20154
rect 2919 20102 2965 20154
rect 2669 20100 2725 20102
rect 2749 20100 2805 20102
rect 2829 20100 2885 20102
rect 2909 20100 2965 20102
rect 2669 19066 2725 19068
rect 2749 19066 2805 19068
rect 2829 19066 2885 19068
rect 2909 19066 2965 19068
rect 2669 19014 2715 19066
rect 2715 19014 2725 19066
rect 2749 19014 2779 19066
rect 2779 19014 2791 19066
rect 2791 19014 2805 19066
rect 2829 19014 2843 19066
rect 2843 19014 2855 19066
rect 2855 19014 2885 19066
rect 2909 19014 2919 19066
rect 2919 19014 2965 19066
rect 2669 19012 2725 19014
rect 2749 19012 2805 19014
rect 2829 19012 2885 19014
rect 2909 19012 2965 19014
rect 2669 17978 2725 17980
rect 2749 17978 2805 17980
rect 2829 17978 2885 17980
rect 2909 17978 2965 17980
rect 2669 17926 2715 17978
rect 2715 17926 2725 17978
rect 2749 17926 2779 17978
rect 2779 17926 2791 17978
rect 2791 17926 2805 17978
rect 2829 17926 2843 17978
rect 2843 17926 2855 17978
rect 2855 17926 2885 17978
rect 2909 17926 2919 17978
rect 2919 17926 2965 17978
rect 2669 17924 2725 17926
rect 2749 17924 2805 17926
rect 2829 17924 2885 17926
rect 2909 17924 2965 17926
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 1858 9424 1914 9480
rect 846 7384 902 7440
rect 1674 8200 1730 8256
rect 846 6604 848 6624
rect 848 6604 900 6624
rect 900 6604 902 6624
rect 846 6568 902 6604
rect 846 5752 902 5808
rect 846 4972 848 4992
rect 848 4972 900 4992
rect 900 4972 902 4992
rect 846 4936 902 4972
rect 754 4120 810 4176
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 12438 42644 12440 42664
rect 12440 42644 12492 42664
rect 12492 42644 12494 42664
rect 3514 18808 3570 18864
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 2502 5616 2558 5672
rect 4382 42458 4438 42460
rect 4462 42458 4518 42460
rect 4542 42458 4598 42460
rect 4622 42458 4678 42460
rect 4382 42406 4428 42458
rect 4428 42406 4438 42458
rect 4462 42406 4492 42458
rect 4492 42406 4504 42458
rect 4504 42406 4518 42458
rect 4542 42406 4556 42458
rect 4556 42406 4568 42458
rect 4568 42406 4598 42458
rect 4622 42406 4632 42458
rect 4632 42406 4678 42458
rect 4382 42404 4438 42406
rect 4462 42404 4518 42406
rect 4542 42404 4598 42406
rect 4622 42404 4678 42406
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 4250 41520 4306 41576
rect 4382 41370 4438 41372
rect 4462 41370 4518 41372
rect 4542 41370 4598 41372
rect 4622 41370 4678 41372
rect 4382 41318 4428 41370
rect 4428 41318 4438 41370
rect 4462 41318 4492 41370
rect 4492 41318 4504 41370
rect 4504 41318 4518 41370
rect 4542 41318 4556 41370
rect 4556 41318 4568 41370
rect 4568 41318 4598 41370
rect 4622 41318 4632 41370
rect 4632 41318 4678 41370
rect 4382 41316 4438 41318
rect 4462 41316 4518 41318
rect 4542 41316 4598 41318
rect 4622 41316 4678 41318
rect 4382 40282 4438 40284
rect 4462 40282 4518 40284
rect 4542 40282 4598 40284
rect 4622 40282 4678 40284
rect 4382 40230 4428 40282
rect 4428 40230 4438 40282
rect 4462 40230 4492 40282
rect 4492 40230 4504 40282
rect 4504 40230 4518 40282
rect 4542 40230 4556 40282
rect 4556 40230 4568 40282
rect 4568 40230 4598 40282
rect 4622 40230 4632 40282
rect 4632 40230 4678 40282
rect 4382 40228 4438 40230
rect 4462 40228 4518 40230
rect 4542 40228 4598 40230
rect 4622 40228 4678 40230
rect 4382 39194 4438 39196
rect 4462 39194 4518 39196
rect 4542 39194 4598 39196
rect 4622 39194 4678 39196
rect 4382 39142 4428 39194
rect 4428 39142 4438 39194
rect 4462 39142 4492 39194
rect 4492 39142 4504 39194
rect 4504 39142 4518 39194
rect 4542 39142 4556 39194
rect 4556 39142 4568 39194
rect 4568 39142 4598 39194
rect 4622 39142 4632 39194
rect 4632 39142 4678 39194
rect 4382 39140 4438 39142
rect 4462 39140 4518 39142
rect 4542 39140 4598 39142
rect 4622 39140 4678 39142
rect 4382 38106 4438 38108
rect 4462 38106 4518 38108
rect 4542 38106 4598 38108
rect 4622 38106 4678 38108
rect 4382 38054 4428 38106
rect 4428 38054 4438 38106
rect 4462 38054 4492 38106
rect 4492 38054 4504 38106
rect 4504 38054 4518 38106
rect 4542 38054 4556 38106
rect 4556 38054 4568 38106
rect 4568 38054 4598 38106
rect 4622 38054 4632 38106
rect 4632 38054 4678 38106
rect 4382 38052 4438 38054
rect 4462 38052 4518 38054
rect 4542 38052 4598 38054
rect 4622 38052 4678 38054
rect 4382 37018 4438 37020
rect 4462 37018 4518 37020
rect 4542 37018 4598 37020
rect 4622 37018 4678 37020
rect 4382 36966 4428 37018
rect 4428 36966 4438 37018
rect 4462 36966 4492 37018
rect 4492 36966 4504 37018
rect 4504 36966 4518 37018
rect 4542 36966 4556 37018
rect 4556 36966 4568 37018
rect 4568 36966 4598 37018
rect 4622 36966 4632 37018
rect 4632 36966 4678 37018
rect 4382 36964 4438 36966
rect 4462 36964 4518 36966
rect 4542 36964 4598 36966
rect 4622 36964 4678 36966
rect 4382 35930 4438 35932
rect 4462 35930 4518 35932
rect 4542 35930 4598 35932
rect 4622 35930 4678 35932
rect 4382 35878 4428 35930
rect 4428 35878 4438 35930
rect 4462 35878 4492 35930
rect 4492 35878 4504 35930
rect 4504 35878 4518 35930
rect 4542 35878 4556 35930
rect 4556 35878 4568 35930
rect 4568 35878 4598 35930
rect 4622 35878 4632 35930
rect 4632 35878 4678 35930
rect 4382 35876 4438 35878
rect 4462 35876 4518 35878
rect 4542 35876 4598 35878
rect 4622 35876 4678 35878
rect 4382 34842 4438 34844
rect 4462 34842 4518 34844
rect 4542 34842 4598 34844
rect 4622 34842 4678 34844
rect 4382 34790 4428 34842
rect 4428 34790 4438 34842
rect 4462 34790 4492 34842
rect 4492 34790 4504 34842
rect 4504 34790 4518 34842
rect 4542 34790 4556 34842
rect 4556 34790 4568 34842
rect 4568 34790 4598 34842
rect 4622 34790 4632 34842
rect 4632 34790 4678 34842
rect 4382 34788 4438 34790
rect 4462 34788 4518 34790
rect 4542 34788 4598 34790
rect 4622 34788 4678 34790
rect 4382 33754 4438 33756
rect 4462 33754 4518 33756
rect 4542 33754 4598 33756
rect 4622 33754 4678 33756
rect 4382 33702 4428 33754
rect 4428 33702 4438 33754
rect 4462 33702 4492 33754
rect 4492 33702 4504 33754
rect 4504 33702 4518 33754
rect 4542 33702 4556 33754
rect 4556 33702 4568 33754
rect 4568 33702 4598 33754
rect 4622 33702 4632 33754
rect 4632 33702 4678 33754
rect 4382 33700 4438 33702
rect 4462 33700 4518 33702
rect 4542 33700 4598 33702
rect 4622 33700 4678 33702
rect 4382 32666 4438 32668
rect 4462 32666 4518 32668
rect 4542 32666 4598 32668
rect 4622 32666 4678 32668
rect 4382 32614 4428 32666
rect 4428 32614 4438 32666
rect 4462 32614 4492 32666
rect 4492 32614 4504 32666
rect 4504 32614 4518 32666
rect 4542 32614 4556 32666
rect 4556 32614 4568 32666
rect 4568 32614 4598 32666
rect 4622 32614 4632 32666
rect 4632 32614 4678 32666
rect 4382 32612 4438 32614
rect 4462 32612 4518 32614
rect 4542 32612 4598 32614
rect 4622 32612 4678 32614
rect 4382 31578 4438 31580
rect 4462 31578 4518 31580
rect 4542 31578 4598 31580
rect 4622 31578 4678 31580
rect 4382 31526 4428 31578
rect 4428 31526 4438 31578
rect 4462 31526 4492 31578
rect 4492 31526 4504 31578
rect 4504 31526 4518 31578
rect 4542 31526 4556 31578
rect 4556 31526 4568 31578
rect 4568 31526 4598 31578
rect 4622 31526 4632 31578
rect 4632 31526 4678 31578
rect 4382 31524 4438 31526
rect 4462 31524 4518 31526
rect 4542 31524 4598 31526
rect 4622 31524 4678 31526
rect 4382 30490 4438 30492
rect 4462 30490 4518 30492
rect 4542 30490 4598 30492
rect 4622 30490 4678 30492
rect 4382 30438 4428 30490
rect 4428 30438 4438 30490
rect 4462 30438 4492 30490
rect 4492 30438 4504 30490
rect 4504 30438 4518 30490
rect 4542 30438 4556 30490
rect 4556 30438 4568 30490
rect 4568 30438 4598 30490
rect 4622 30438 4632 30490
rect 4632 30438 4678 30490
rect 4382 30436 4438 30438
rect 4462 30436 4518 30438
rect 4542 30436 4598 30438
rect 4622 30436 4678 30438
rect 4382 29402 4438 29404
rect 4462 29402 4518 29404
rect 4542 29402 4598 29404
rect 4622 29402 4678 29404
rect 4382 29350 4428 29402
rect 4428 29350 4438 29402
rect 4462 29350 4492 29402
rect 4492 29350 4504 29402
rect 4504 29350 4518 29402
rect 4542 29350 4556 29402
rect 4556 29350 4568 29402
rect 4568 29350 4598 29402
rect 4622 29350 4632 29402
rect 4632 29350 4678 29402
rect 4382 29348 4438 29350
rect 4462 29348 4518 29350
rect 4542 29348 4598 29350
rect 4622 29348 4678 29350
rect 4382 28314 4438 28316
rect 4462 28314 4518 28316
rect 4542 28314 4598 28316
rect 4622 28314 4678 28316
rect 4382 28262 4428 28314
rect 4428 28262 4438 28314
rect 4462 28262 4492 28314
rect 4492 28262 4504 28314
rect 4504 28262 4518 28314
rect 4542 28262 4556 28314
rect 4556 28262 4568 28314
rect 4568 28262 4598 28314
rect 4622 28262 4632 28314
rect 4632 28262 4678 28314
rect 4382 28260 4438 28262
rect 4462 28260 4518 28262
rect 4542 28260 4598 28262
rect 4622 28260 4678 28262
rect 4382 27226 4438 27228
rect 4462 27226 4518 27228
rect 4542 27226 4598 27228
rect 4622 27226 4678 27228
rect 4382 27174 4428 27226
rect 4428 27174 4438 27226
rect 4462 27174 4492 27226
rect 4492 27174 4504 27226
rect 4504 27174 4518 27226
rect 4542 27174 4556 27226
rect 4556 27174 4568 27226
rect 4568 27174 4598 27226
rect 4622 27174 4632 27226
rect 4632 27174 4678 27226
rect 4382 27172 4438 27174
rect 4462 27172 4518 27174
rect 4542 27172 4598 27174
rect 4622 27172 4678 27174
rect 4382 26138 4438 26140
rect 4462 26138 4518 26140
rect 4542 26138 4598 26140
rect 4622 26138 4678 26140
rect 4382 26086 4428 26138
rect 4428 26086 4438 26138
rect 4462 26086 4492 26138
rect 4492 26086 4504 26138
rect 4504 26086 4518 26138
rect 4542 26086 4556 26138
rect 4556 26086 4568 26138
rect 4568 26086 4598 26138
rect 4622 26086 4632 26138
rect 4632 26086 4678 26138
rect 4382 26084 4438 26086
rect 4462 26084 4518 26086
rect 4542 26084 4598 26086
rect 4622 26084 4678 26086
rect 4382 25050 4438 25052
rect 4462 25050 4518 25052
rect 4542 25050 4598 25052
rect 4622 25050 4678 25052
rect 4382 24998 4428 25050
rect 4428 24998 4438 25050
rect 4462 24998 4492 25050
rect 4492 24998 4504 25050
rect 4504 24998 4518 25050
rect 4542 24998 4556 25050
rect 4556 24998 4568 25050
rect 4568 24998 4598 25050
rect 4622 24998 4632 25050
rect 4632 24998 4678 25050
rect 4382 24996 4438 24998
rect 4462 24996 4518 24998
rect 4542 24996 4598 24998
rect 4622 24996 4678 24998
rect 4382 23962 4438 23964
rect 4462 23962 4518 23964
rect 4542 23962 4598 23964
rect 4622 23962 4678 23964
rect 4382 23910 4428 23962
rect 4428 23910 4438 23962
rect 4462 23910 4492 23962
rect 4492 23910 4504 23962
rect 4504 23910 4518 23962
rect 4542 23910 4556 23962
rect 4556 23910 4568 23962
rect 4568 23910 4598 23962
rect 4622 23910 4632 23962
rect 4632 23910 4678 23962
rect 4382 23908 4438 23910
rect 4462 23908 4518 23910
rect 4542 23908 4598 23910
rect 4622 23908 4678 23910
rect 4382 22874 4438 22876
rect 4462 22874 4518 22876
rect 4542 22874 4598 22876
rect 4622 22874 4678 22876
rect 4382 22822 4428 22874
rect 4428 22822 4438 22874
rect 4462 22822 4492 22874
rect 4492 22822 4504 22874
rect 4504 22822 4518 22874
rect 4542 22822 4556 22874
rect 4556 22822 4568 22874
rect 4568 22822 4598 22874
rect 4622 22822 4632 22874
rect 4632 22822 4678 22874
rect 4382 22820 4438 22822
rect 4462 22820 4518 22822
rect 4542 22820 4598 22822
rect 4622 22820 4678 22822
rect 4382 21786 4438 21788
rect 4462 21786 4518 21788
rect 4542 21786 4598 21788
rect 4622 21786 4678 21788
rect 4382 21734 4428 21786
rect 4428 21734 4438 21786
rect 4462 21734 4492 21786
rect 4492 21734 4504 21786
rect 4504 21734 4518 21786
rect 4542 21734 4556 21786
rect 4556 21734 4568 21786
rect 4568 21734 4598 21786
rect 4622 21734 4632 21786
rect 4632 21734 4678 21786
rect 4382 21732 4438 21734
rect 4462 21732 4518 21734
rect 4542 21732 4598 21734
rect 4622 21732 4678 21734
rect 4382 20698 4438 20700
rect 4462 20698 4518 20700
rect 4542 20698 4598 20700
rect 4622 20698 4678 20700
rect 4382 20646 4428 20698
rect 4428 20646 4438 20698
rect 4462 20646 4492 20698
rect 4492 20646 4504 20698
rect 4504 20646 4518 20698
rect 4542 20646 4556 20698
rect 4556 20646 4568 20698
rect 4568 20646 4598 20698
rect 4622 20646 4632 20698
rect 4632 20646 4678 20698
rect 4382 20644 4438 20646
rect 4462 20644 4518 20646
rect 4542 20644 4598 20646
rect 4622 20644 4678 20646
rect 7809 42458 7865 42460
rect 7889 42458 7945 42460
rect 7969 42458 8025 42460
rect 8049 42458 8105 42460
rect 7809 42406 7855 42458
rect 7855 42406 7865 42458
rect 7889 42406 7919 42458
rect 7919 42406 7931 42458
rect 7931 42406 7945 42458
rect 7969 42406 7983 42458
rect 7983 42406 7995 42458
rect 7995 42406 8025 42458
rect 8049 42406 8059 42458
rect 8059 42406 8105 42458
rect 7809 42404 7865 42406
rect 7889 42404 7945 42406
rect 7969 42404 8025 42406
rect 8049 42404 8105 42406
rect 6096 41914 6152 41916
rect 6176 41914 6232 41916
rect 6256 41914 6312 41916
rect 6336 41914 6392 41916
rect 6096 41862 6142 41914
rect 6142 41862 6152 41914
rect 6176 41862 6206 41914
rect 6206 41862 6218 41914
rect 6218 41862 6232 41914
rect 6256 41862 6270 41914
rect 6270 41862 6282 41914
rect 6282 41862 6312 41914
rect 6336 41862 6346 41914
rect 6346 41862 6392 41914
rect 6096 41860 6152 41862
rect 6176 41860 6232 41862
rect 6256 41860 6312 41862
rect 6336 41860 6392 41862
rect 9523 41914 9579 41916
rect 9603 41914 9659 41916
rect 9683 41914 9739 41916
rect 9763 41914 9819 41916
rect 9523 41862 9569 41914
rect 9569 41862 9579 41914
rect 9603 41862 9633 41914
rect 9633 41862 9645 41914
rect 9645 41862 9659 41914
rect 9683 41862 9697 41914
rect 9697 41862 9709 41914
rect 9709 41862 9739 41914
rect 9763 41862 9773 41914
rect 9773 41862 9819 41914
rect 9523 41860 9579 41862
rect 9603 41860 9659 41862
rect 9683 41860 9739 41862
rect 9763 41860 9819 41862
rect 9402 41656 9458 41712
rect 11236 42458 11292 42460
rect 11316 42458 11372 42460
rect 11396 42458 11452 42460
rect 11476 42458 11532 42460
rect 11236 42406 11282 42458
rect 11282 42406 11292 42458
rect 11316 42406 11346 42458
rect 11346 42406 11358 42458
rect 11358 42406 11372 42458
rect 11396 42406 11410 42458
rect 11410 42406 11422 42458
rect 11422 42406 11452 42458
rect 11476 42406 11486 42458
rect 11486 42406 11532 42458
rect 11236 42404 11292 42406
rect 11316 42404 11372 42406
rect 11396 42404 11452 42406
rect 11476 42404 11532 42406
rect 12438 42608 12494 42644
rect 14663 43546 14719 43548
rect 14743 43546 14799 43548
rect 14823 43546 14879 43548
rect 14903 43546 14959 43548
rect 14663 43494 14709 43546
rect 14709 43494 14719 43546
rect 14743 43494 14773 43546
rect 14773 43494 14785 43546
rect 14785 43494 14799 43546
rect 14823 43494 14837 43546
rect 14837 43494 14849 43546
rect 14849 43494 14879 43546
rect 14903 43494 14913 43546
rect 14913 43494 14959 43546
rect 14663 43492 14719 43494
rect 14743 43492 14799 43494
rect 14823 43492 14879 43494
rect 14903 43492 14959 43494
rect 14663 42458 14719 42460
rect 14743 42458 14799 42460
rect 14823 42458 14879 42460
rect 14903 42458 14959 42460
rect 14663 42406 14709 42458
rect 14709 42406 14719 42458
rect 14743 42406 14773 42458
rect 14773 42406 14785 42458
rect 14785 42406 14799 42458
rect 14823 42406 14837 42458
rect 14837 42406 14849 42458
rect 14849 42406 14879 42458
rect 14903 42406 14913 42458
rect 14913 42406 14959 42458
rect 14663 42404 14719 42406
rect 14743 42404 14799 42406
rect 14823 42404 14879 42406
rect 14903 42404 14959 42406
rect 12950 41914 13006 41916
rect 13030 41914 13086 41916
rect 13110 41914 13166 41916
rect 13190 41914 13246 41916
rect 12950 41862 12996 41914
rect 12996 41862 13006 41914
rect 13030 41862 13060 41914
rect 13060 41862 13072 41914
rect 13072 41862 13086 41914
rect 13110 41862 13124 41914
rect 13124 41862 13136 41914
rect 13136 41862 13166 41914
rect 13190 41862 13200 41914
rect 13200 41862 13246 41914
rect 12950 41860 13006 41862
rect 13030 41860 13086 41862
rect 13110 41860 13166 41862
rect 13190 41860 13246 41862
rect 11702 41520 11758 41576
rect 5078 41384 5134 41440
rect 10966 41384 11022 41440
rect 7809 41370 7865 41372
rect 7889 41370 7945 41372
rect 7969 41370 8025 41372
rect 8049 41370 8105 41372
rect 7809 41318 7855 41370
rect 7855 41318 7865 41370
rect 7889 41318 7919 41370
rect 7919 41318 7931 41370
rect 7931 41318 7945 41370
rect 7969 41318 7983 41370
rect 7983 41318 7995 41370
rect 7995 41318 8025 41370
rect 8049 41318 8059 41370
rect 8059 41318 8105 41370
rect 7809 41316 7865 41318
rect 7889 41316 7945 41318
rect 7969 41316 8025 41318
rect 8049 41316 8105 41318
rect 11236 41370 11292 41372
rect 11316 41370 11372 41372
rect 11396 41370 11452 41372
rect 11476 41370 11532 41372
rect 11236 41318 11282 41370
rect 11282 41318 11292 41370
rect 11316 41318 11346 41370
rect 11346 41318 11358 41370
rect 11358 41318 11372 41370
rect 11396 41318 11410 41370
rect 11410 41318 11422 41370
rect 11422 41318 11452 41370
rect 11476 41318 11486 41370
rect 11486 41318 11532 41370
rect 11236 41316 11292 41318
rect 11316 41316 11372 41318
rect 11396 41316 11452 41318
rect 11476 41316 11532 41318
rect 6096 40826 6152 40828
rect 6176 40826 6232 40828
rect 6256 40826 6312 40828
rect 6336 40826 6392 40828
rect 6096 40774 6142 40826
rect 6142 40774 6152 40826
rect 6176 40774 6206 40826
rect 6206 40774 6218 40826
rect 6218 40774 6232 40826
rect 6256 40774 6270 40826
rect 6270 40774 6282 40826
rect 6282 40774 6312 40826
rect 6336 40774 6346 40826
rect 6346 40774 6392 40826
rect 6096 40772 6152 40774
rect 6176 40772 6232 40774
rect 6256 40772 6312 40774
rect 6336 40772 6392 40774
rect 7809 40282 7865 40284
rect 7889 40282 7945 40284
rect 7969 40282 8025 40284
rect 8049 40282 8105 40284
rect 7809 40230 7855 40282
rect 7855 40230 7865 40282
rect 7889 40230 7919 40282
rect 7919 40230 7931 40282
rect 7931 40230 7945 40282
rect 7969 40230 7983 40282
rect 7983 40230 7995 40282
rect 7995 40230 8025 40282
rect 8049 40230 8059 40282
rect 8059 40230 8105 40282
rect 7809 40228 7865 40230
rect 7889 40228 7945 40230
rect 7969 40228 8025 40230
rect 8049 40228 8105 40230
rect 9523 40826 9579 40828
rect 9603 40826 9659 40828
rect 9683 40826 9739 40828
rect 9763 40826 9819 40828
rect 9523 40774 9569 40826
rect 9569 40774 9579 40826
rect 9603 40774 9633 40826
rect 9633 40774 9645 40826
rect 9645 40774 9659 40826
rect 9683 40774 9697 40826
rect 9697 40774 9709 40826
rect 9709 40774 9739 40826
rect 9763 40774 9773 40826
rect 9773 40774 9819 40826
rect 9523 40772 9579 40774
rect 9603 40772 9659 40774
rect 9683 40772 9739 40774
rect 9763 40772 9819 40774
rect 12950 40826 13006 40828
rect 13030 40826 13086 40828
rect 13110 40826 13166 40828
rect 13190 40826 13246 40828
rect 12950 40774 12996 40826
rect 12996 40774 13006 40826
rect 13030 40774 13060 40826
rect 13060 40774 13072 40826
rect 13072 40774 13086 40826
rect 13110 40774 13124 40826
rect 13124 40774 13136 40826
rect 13136 40774 13166 40826
rect 13190 40774 13200 40826
rect 13200 40774 13246 40826
rect 12950 40772 13006 40774
rect 13030 40772 13086 40774
rect 13110 40772 13166 40774
rect 13190 40772 13246 40774
rect 11236 40282 11292 40284
rect 11316 40282 11372 40284
rect 11396 40282 11452 40284
rect 11476 40282 11532 40284
rect 11236 40230 11282 40282
rect 11282 40230 11292 40282
rect 11316 40230 11346 40282
rect 11346 40230 11358 40282
rect 11358 40230 11372 40282
rect 11396 40230 11410 40282
rect 11410 40230 11422 40282
rect 11422 40230 11452 40282
rect 11476 40230 11486 40282
rect 11486 40230 11532 40282
rect 11236 40228 11292 40230
rect 11316 40228 11372 40230
rect 11396 40228 11452 40230
rect 11476 40228 11532 40230
rect 9310 40044 9366 40080
rect 9310 40024 9312 40044
rect 9312 40024 9364 40044
rect 9364 40024 9366 40044
rect 6096 39738 6152 39740
rect 6176 39738 6232 39740
rect 6256 39738 6312 39740
rect 6336 39738 6392 39740
rect 6096 39686 6142 39738
rect 6142 39686 6152 39738
rect 6176 39686 6206 39738
rect 6206 39686 6218 39738
rect 6218 39686 6232 39738
rect 6256 39686 6270 39738
rect 6270 39686 6282 39738
rect 6282 39686 6312 39738
rect 6336 39686 6346 39738
rect 6346 39686 6392 39738
rect 6096 39684 6152 39686
rect 6176 39684 6232 39686
rect 6256 39684 6312 39686
rect 6336 39684 6392 39686
rect 9523 39738 9579 39740
rect 9603 39738 9659 39740
rect 9683 39738 9739 39740
rect 9763 39738 9819 39740
rect 9523 39686 9569 39738
rect 9569 39686 9579 39738
rect 9603 39686 9633 39738
rect 9633 39686 9645 39738
rect 9645 39686 9659 39738
rect 9683 39686 9697 39738
rect 9697 39686 9709 39738
rect 9709 39686 9739 39738
rect 9763 39686 9773 39738
rect 9773 39686 9819 39738
rect 9523 39684 9579 39686
rect 9603 39684 9659 39686
rect 9683 39684 9739 39686
rect 9763 39684 9819 39686
rect 12950 39738 13006 39740
rect 13030 39738 13086 39740
rect 13110 39738 13166 39740
rect 13190 39738 13246 39740
rect 12950 39686 12996 39738
rect 12996 39686 13006 39738
rect 13030 39686 13060 39738
rect 13060 39686 13072 39738
rect 13072 39686 13086 39738
rect 13110 39686 13124 39738
rect 13124 39686 13136 39738
rect 13136 39686 13166 39738
rect 13190 39686 13200 39738
rect 13200 39686 13246 39738
rect 12950 39684 13006 39686
rect 13030 39684 13086 39686
rect 13110 39684 13166 39686
rect 13190 39684 13246 39686
rect 13726 39752 13782 39808
rect 14002 39480 14058 39536
rect 14186 39480 14242 39536
rect 4382 19610 4438 19612
rect 4462 19610 4518 19612
rect 4542 19610 4598 19612
rect 4622 19610 4678 19612
rect 4382 19558 4428 19610
rect 4428 19558 4438 19610
rect 4462 19558 4492 19610
rect 4492 19558 4504 19610
rect 4504 19558 4518 19610
rect 4542 19558 4556 19610
rect 4556 19558 4568 19610
rect 4568 19558 4598 19610
rect 4622 19558 4632 19610
rect 4632 19558 4678 19610
rect 4382 19556 4438 19558
rect 4462 19556 4518 19558
rect 4542 19556 4598 19558
rect 4622 19556 4678 19558
rect 4382 18522 4438 18524
rect 4462 18522 4518 18524
rect 4542 18522 4598 18524
rect 4622 18522 4678 18524
rect 4382 18470 4428 18522
rect 4428 18470 4438 18522
rect 4462 18470 4492 18522
rect 4492 18470 4504 18522
rect 4504 18470 4518 18522
rect 4542 18470 4556 18522
rect 4556 18470 4568 18522
rect 4568 18470 4598 18522
rect 4622 18470 4632 18522
rect 4632 18470 4678 18522
rect 4382 18468 4438 18470
rect 4462 18468 4518 18470
rect 4542 18468 4598 18470
rect 4622 18468 4678 18470
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 7809 39194 7865 39196
rect 7889 39194 7945 39196
rect 7969 39194 8025 39196
rect 8049 39194 8105 39196
rect 7809 39142 7855 39194
rect 7855 39142 7865 39194
rect 7889 39142 7919 39194
rect 7919 39142 7931 39194
rect 7931 39142 7945 39194
rect 7969 39142 7983 39194
rect 7983 39142 7995 39194
rect 7995 39142 8025 39194
rect 8049 39142 8059 39194
rect 8059 39142 8105 39194
rect 7809 39140 7865 39142
rect 7889 39140 7945 39142
rect 7969 39140 8025 39142
rect 8049 39140 8105 39142
rect 11236 39194 11292 39196
rect 11316 39194 11372 39196
rect 11396 39194 11452 39196
rect 11476 39194 11532 39196
rect 11236 39142 11282 39194
rect 11282 39142 11292 39194
rect 11316 39142 11346 39194
rect 11346 39142 11358 39194
rect 11358 39142 11372 39194
rect 11396 39142 11410 39194
rect 11410 39142 11422 39194
rect 11422 39142 11452 39194
rect 11476 39142 11486 39194
rect 11486 39142 11532 39194
rect 11236 39140 11292 39142
rect 11316 39140 11372 39142
rect 11396 39140 11452 39142
rect 11476 39140 11532 39142
rect 6096 38650 6152 38652
rect 6176 38650 6232 38652
rect 6256 38650 6312 38652
rect 6336 38650 6392 38652
rect 6096 38598 6142 38650
rect 6142 38598 6152 38650
rect 6176 38598 6206 38650
rect 6206 38598 6218 38650
rect 6218 38598 6232 38650
rect 6256 38598 6270 38650
rect 6270 38598 6282 38650
rect 6282 38598 6312 38650
rect 6336 38598 6346 38650
rect 6346 38598 6392 38650
rect 6096 38596 6152 38598
rect 6176 38596 6232 38598
rect 6256 38596 6312 38598
rect 6336 38596 6392 38598
rect 9523 38650 9579 38652
rect 9603 38650 9659 38652
rect 9683 38650 9739 38652
rect 9763 38650 9819 38652
rect 9523 38598 9569 38650
rect 9569 38598 9579 38650
rect 9603 38598 9633 38650
rect 9633 38598 9645 38650
rect 9645 38598 9659 38650
rect 9683 38598 9697 38650
rect 9697 38598 9709 38650
rect 9709 38598 9739 38650
rect 9763 38598 9773 38650
rect 9773 38598 9819 38650
rect 9523 38596 9579 38598
rect 9603 38596 9659 38598
rect 9683 38596 9739 38598
rect 9763 38596 9819 38598
rect 7809 38106 7865 38108
rect 7889 38106 7945 38108
rect 7969 38106 8025 38108
rect 8049 38106 8105 38108
rect 7809 38054 7855 38106
rect 7855 38054 7865 38106
rect 7889 38054 7919 38106
rect 7919 38054 7931 38106
rect 7931 38054 7945 38106
rect 7969 38054 7983 38106
rect 7983 38054 7995 38106
rect 7995 38054 8025 38106
rect 8049 38054 8059 38106
rect 8059 38054 8105 38106
rect 7809 38052 7865 38054
rect 7889 38052 7945 38054
rect 7969 38052 8025 38054
rect 8049 38052 8105 38054
rect 11236 38106 11292 38108
rect 11316 38106 11372 38108
rect 11396 38106 11452 38108
rect 11476 38106 11532 38108
rect 11236 38054 11282 38106
rect 11282 38054 11292 38106
rect 11316 38054 11346 38106
rect 11346 38054 11358 38106
rect 11358 38054 11372 38106
rect 11396 38054 11410 38106
rect 11410 38054 11422 38106
rect 11422 38054 11452 38106
rect 11476 38054 11486 38106
rect 11486 38054 11532 38106
rect 11236 38052 11292 38054
rect 11316 38052 11372 38054
rect 11396 38052 11452 38054
rect 11476 38052 11532 38054
rect 6096 37562 6152 37564
rect 6176 37562 6232 37564
rect 6256 37562 6312 37564
rect 6336 37562 6392 37564
rect 6096 37510 6142 37562
rect 6142 37510 6152 37562
rect 6176 37510 6206 37562
rect 6206 37510 6218 37562
rect 6218 37510 6232 37562
rect 6256 37510 6270 37562
rect 6270 37510 6282 37562
rect 6282 37510 6312 37562
rect 6336 37510 6346 37562
rect 6346 37510 6392 37562
rect 6096 37508 6152 37510
rect 6176 37508 6232 37510
rect 6256 37508 6312 37510
rect 6336 37508 6392 37510
rect 6826 36624 6882 36680
rect 6096 36474 6152 36476
rect 6176 36474 6232 36476
rect 6256 36474 6312 36476
rect 6336 36474 6392 36476
rect 6096 36422 6142 36474
rect 6142 36422 6152 36474
rect 6176 36422 6206 36474
rect 6206 36422 6218 36474
rect 6218 36422 6232 36474
rect 6256 36422 6270 36474
rect 6270 36422 6282 36474
rect 6282 36422 6312 36474
rect 6336 36422 6346 36474
rect 6346 36422 6392 36474
rect 6096 36420 6152 36422
rect 6176 36420 6232 36422
rect 6256 36420 6312 36422
rect 6336 36420 6392 36422
rect 5630 29144 5686 29200
rect 6096 35386 6152 35388
rect 6176 35386 6232 35388
rect 6256 35386 6312 35388
rect 6336 35386 6392 35388
rect 6096 35334 6142 35386
rect 6142 35334 6152 35386
rect 6176 35334 6206 35386
rect 6206 35334 6218 35386
rect 6218 35334 6232 35386
rect 6256 35334 6270 35386
rect 6270 35334 6282 35386
rect 6282 35334 6312 35386
rect 6336 35334 6346 35386
rect 6346 35334 6392 35386
rect 6096 35332 6152 35334
rect 6176 35332 6232 35334
rect 6256 35332 6312 35334
rect 6336 35332 6392 35334
rect 5998 35128 6054 35184
rect 6096 34298 6152 34300
rect 6176 34298 6232 34300
rect 6256 34298 6312 34300
rect 6336 34298 6392 34300
rect 6096 34246 6142 34298
rect 6142 34246 6152 34298
rect 6176 34246 6206 34298
rect 6206 34246 6218 34298
rect 6218 34246 6232 34298
rect 6256 34246 6270 34298
rect 6270 34246 6282 34298
rect 6282 34246 6312 34298
rect 6336 34246 6346 34298
rect 6346 34246 6392 34298
rect 6096 34244 6152 34246
rect 6176 34244 6232 34246
rect 6256 34244 6312 34246
rect 6336 34244 6392 34246
rect 6096 33210 6152 33212
rect 6176 33210 6232 33212
rect 6256 33210 6312 33212
rect 6336 33210 6392 33212
rect 6096 33158 6142 33210
rect 6142 33158 6152 33210
rect 6176 33158 6206 33210
rect 6206 33158 6218 33210
rect 6218 33158 6232 33210
rect 6256 33158 6270 33210
rect 6270 33158 6282 33210
rect 6282 33158 6312 33210
rect 6336 33158 6346 33210
rect 6346 33158 6392 33210
rect 6096 33156 6152 33158
rect 6176 33156 6232 33158
rect 6256 33156 6312 33158
rect 6336 33156 6392 33158
rect 6096 32122 6152 32124
rect 6176 32122 6232 32124
rect 6256 32122 6312 32124
rect 6336 32122 6392 32124
rect 6096 32070 6142 32122
rect 6142 32070 6152 32122
rect 6176 32070 6206 32122
rect 6206 32070 6218 32122
rect 6218 32070 6232 32122
rect 6256 32070 6270 32122
rect 6270 32070 6282 32122
rect 6282 32070 6312 32122
rect 6336 32070 6346 32122
rect 6346 32070 6392 32122
rect 6096 32068 6152 32070
rect 6176 32068 6232 32070
rect 6256 32068 6312 32070
rect 6336 32068 6392 32070
rect 6918 32272 6974 32328
rect 6096 31034 6152 31036
rect 6176 31034 6232 31036
rect 6256 31034 6312 31036
rect 6336 31034 6392 31036
rect 6096 30982 6142 31034
rect 6142 30982 6152 31034
rect 6176 30982 6206 31034
rect 6206 30982 6218 31034
rect 6218 30982 6232 31034
rect 6256 30982 6270 31034
rect 6270 30982 6282 31034
rect 6282 30982 6312 31034
rect 6336 30982 6346 31034
rect 6346 30982 6392 31034
rect 6096 30980 6152 30982
rect 6176 30980 6232 30982
rect 6256 30980 6312 30982
rect 6336 30980 6392 30982
rect 6096 29946 6152 29948
rect 6176 29946 6232 29948
rect 6256 29946 6312 29948
rect 6336 29946 6392 29948
rect 6096 29894 6142 29946
rect 6142 29894 6152 29946
rect 6176 29894 6206 29946
rect 6206 29894 6218 29946
rect 6218 29894 6232 29946
rect 6256 29894 6270 29946
rect 6270 29894 6282 29946
rect 6282 29894 6312 29946
rect 6336 29894 6346 29946
rect 6346 29894 6392 29946
rect 6096 29892 6152 29894
rect 6176 29892 6232 29894
rect 6256 29892 6312 29894
rect 6336 29892 6392 29894
rect 6096 28858 6152 28860
rect 6176 28858 6232 28860
rect 6256 28858 6312 28860
rect 6336 28858 6392 28860
rect 6096 28806 6142 28858
rect 6142 28806 6152 28858
rect 6176 28806 6206 28858
rect 6206 28806 6218 28858
rect 6218 28806 6232 28858
rect 6256 28806 6270 28858
rect 6270 28806 6282 28858
rect 6282 28806 6312 28858
rect 6336 28806 6346 28858
rect 6346 28806 6392 28858
rect 6096 28804 6152 28806
rect 6176 28804 6232 28806
rect 6256 28804 6312 28806
rect 6336 28804 6392 28806
rect 6096 27770 6152 27772
rect 6176 27770 6232 27772
rect 6256 27770 6312 27772
rect 6336 27770 6392 27772
rect 6096 27718 6142 27770
rect 6142 27718 6152 27770
rect 6176 27718 6206 27770
rect 6206 27718 6218 27770
rect 6218 27718 6232 27770
rect 6256 27718 6270 27770
rect 6270 27718 6282 27770
rect 6282 27718 6312 27770
rect 6336 27718 6346 27770
rect 6346 27718 6392 27770
rect 6096 27716 6152 27718
rect 6176 27716 6232 27718
rect 6256 27716 6312 27718
rect 6336 27716 6392 27718
rect 6096 26682 6152 26684
rect 6176 26682 6232 26684
rect 6256 26682 6312 26684
rect 6336 26682 6392 26684
rect 6096 26630 6142 26682
rect 6142 26630 6152 26682
rect 6176 26630 6206 26682
rect 6206 26630 6218 26682
rect 6218 26630 6232 26682
rect 6256 26630 6270 26682
rect 6270 26630 6282 26682
rect 6282 26630 6312 26682
rect 6336 26630 6346 26682
rect 6346 26630 6392 26682
rect 6096 26628 6152 26630
rect 6176 26628 6232 26630
rect 6256 26628 6312 26630
rect 6336 26628 6392 26630
rect 6096 25594 6152 25596
rect 6176 25594 6232 25596
rect 6256 25594 6312 25596
rect 6336 25594 6392 25596
rect 6096 25542 6142 25594
rect 6142 25542 6152 25594
rect 6176 25542 6206 25594
rect 6206 25542 6218 25594
rect 6218 25542 6232 25594
rect 6256 25542 6270 25594
rect 6270 25542 6282 25594
rect 6282 25542 6312 25594
rect 6336 25542 6346 25594
rect 6346 25542 6392 25594
rect 6096 25540 6152 25542
rect 6176 25540 6232 25542
rect 6256 25540 6312 25542
rect 6336 25540 6392 25542
rect 5538 19352 5594 19408
rect 6096 24506 6152 24508
rect 6176 24506 6232 24508
rect 6256 24506 6312 24508
rect 6336 24506 6392 24508
rect 6096 24454 6142 24506
rect 6142 24454 6152 24506
rect 6176 24454 6206 24506
rect 6206 24454 6218 24506
rect 6218 24454 6232 24506
rect 6256 24454 6270 24506
rect 6270 24454 6282 24506
rect 6282 24454 6312 24506
rect 6336 24454 6346 24506
rect 6346 24454 6392 24506
rect 6096 24452 6152 24454
rect 6176 24452 6232 24454
rect 6256 24452 6312 24454
rect 6336 24452 6392 24454
rect 5906 24248 5962 24304
rect 5446 17720 5502 17776
rect 5170 17040 5226 17096
rect 5446 8336 5502 8392
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 6096 23418 6152 23420
rect 6176 23418 6232 23420
rect 6256 23418 6312 23420
rect 6336 23418 6392 23420
rect 6096 23366 6142 23418
rect 6142 23366 6152 23418
rect 6176 23366 6206 23418
rect 6206 23366 6218 23418
rect 6218 23366 6232 23418
rect 6256 23366 6270 23418
rect 6270 23366 6282 23418
rect 6282 23366 6312 23418
rect 6336 23366 6346 23418
rect 6346 23366 6392 23418
rect 6096 23364 6152 23366
rect 6176 23364 6232 23366
rect 6256 23364 6312 23366
rect 6336 23364 6392 23366
rect 6096 22330 6152 22332
rect 6176 22330 6232 22332
rect 6256 22330 6312 22332
rect 6336 22330 6392 22332
rect 6096 22278 6142 22330
rect 6142 22278 6152 22330
rect 6176 22278 6206 22330
rect 6206 22278 6218 22330
rect 6218 22278 6232 22330
rect 6256 22278 6270 22330
rect 6270 22278 6282 22330
rect 6282 22278 6312 22330
rect 6336 22278 6346 22330
rect 6346 22278 6392 22330
rect 6096 22276 6152 22278
rect 6176 22276 6232 22278
rect 6256 22276 6312 22278
rect 6336 22276 6392 22278
rect 6274 21528 6330 21584
rect 6096 21242 6152 21244
rect 6176 21242 6232 21244
rect 6256 21242 6312 21244
rect 6336 21242 6392 21244
rect 6096 21190 6142 21242
rect 6142 21190 6152 21242
rect 6176 21190 6206 21242
rect 6206 21190 6218 21242
rect 6218 21190 6232 21242
rect 6256 21190 6270 21242
rect 6270 21190 6282 21242
rect 6282 21190 6312 21242
rect 6336 21190 6346 21242
rect 6346 21190 6392 21242
rect 6096 21188 6152 21190
rect 6176 21188 6232 21190
rect 6256 21188 6312 21190
rect 6336 21188 6392 21190
rect 6096 20154 6152 20156
rect 6176 20154 6232 20156
rect 6256 20154 6312 20156
rect 6336 20154 6392 20156
rect 6096 20102 6142 20154
rect 6142 20102 6152 20154
rect 6176 20102 6206 20154
rect 6206 20102 6218 20154
rect 6218 20102 6232 20154
rect 6256 20102 6270 20154
rect 6270 20102 6282 20154
rect 6282 20102 6312 20154
rect 6336 20102 6346 20154
rect 6346 20102 6392 20154
rect 6096 20100 6152 20102
rect 6176 20100 6232 20102
rect 6256 20100 6312 20102
rect 6336 20100 6392 20102
rect 6096 19066 6152 19068
rect 6176 19066 6232 19068
rect 6256 19066 6312 19068
rect 6336 19066 6392 19068
rect 6096 19014 6142 19066
rect 6142 19014 6152 19066
rect 6176 19014 6206 19066
rect 6206 19014 6218 19066
rect 6218 19014 6232 19066
rect 6256 19014 6270 19066
rect 6270 19014 6282 19066
rect 6282 19014 6312 19066
rect 6336 19014 6346 19066
rect 6346 19014 6392 19066
rect 6096 19012 6152 19014
rect 6176 19012 6232 19014
rect 6256 19012 6312 19014
rect 6336 19012 6392 19014
rect 6096 17978 6152 17980
rect 6176 17978 6232 17980
rect 6256 17978 6312 17980
rect 6336 17978 6392 17980
rect 6096 17926 6142 17978
rect 6142 17926 6152 17978
rect 6176 17926 6206 17978
rect 6206 17926 6218 17978
rect 6218 17926 6232 17978
rect 6256 17926 6270 17978
rect 6270 17926 6282 17978
rect 6282 17926 6312 17978
rect 6336 17926 6346 17978
rect 6346 17926 6392 17978
rect 6096 17924 6152 17926
rect 6176 17924 6232 17926
rect 6256 17924 6312 17926
rect 6336 17924 6392 17926
rect 7194 23976 7250 24032
rect 7102 23840 7158 23896
rect 9523 37562 9579 37564
rect 9603 37562 9659 37564
rect 9683 37562 9739 37564
rect 9763 37562 9819 37564
rect 9523 37510 9569 37562
rect 9569 37510 9579 37562
rect 9603 37510 9633 37562
rect 9633 37510 9645 37562
rect 9645 37510 9659 37562
rect 9683 37510 9697 37562
rect 9697 37510 9709 37562
rect 9709 37510 9739 37562
rect 9763 37510 9773 37562
rect 9773 37510 9819 37562
rect 9523 37508 9579 37510
rect 9603 37508 9659 37510
rect 9683 37508 9739 37510
rect 9763 37508 9819 37510
rect 9862 37168 9918 37224
rect 7809 37018 7865 37020
rect 7889 37018 7945 37020
rect 7969 37018 8025 37020
rect 8049 37018 8105 37020
rect 7809 36966 7855 37018
rect 7855 36966 7865 37018
rect 7889 36966 7919 37018
rect 7919 36966 7931 37018
rect 7931 36966 7945 37018
rect 7969 36966 7983 37018
rect 7983 36966 7995 37018
rect 7995 36966 8025 37018
rect 8049 36966 8059 37018
rect 8059 36966 8105 37018
rect 7809 36964 7865 36966
rect 7889 36964 7945 36966
rect 7969 36964 8025 36966
rect 8049 36964 8105 36966
rect 9523 36474 9579 36476
rect 9603 36474 9659 36476
rect 9683 36474 9739 36476
rect 9763 36474 9819 36476
rect 9523 36422 9569 36474
rect 9569 36422 9579 36474
rect 9603 36422 9633 36474
rect 9633 36422 9645 36474
rect 9645 36422 9659 36474
rect 9683 36422 9697 36474
rect 9697 36422 9709 36474
rect 9709 36422 9739 36474
rect 9763 36422 9773 36474
rect 9773 36422 9819 36474
rect 9523 36420 9579 36422
rect 9603 36420 9659 36422
rect 9683 36420 9739 36422
rect 9763 36420 9819 36422
rect 7809 35930 7865 35932
rect 7889 35930 7945 35932
rect 7969 35930 8025 35932
rect 8049 35930 8105 35932
rect 7809 35878 7855 35930
rect 7855 35878 7865 35930
rect 7889 35878 7919 35930
rect 7919 35878 7931 35930
rect 7931 35878 7945 35930
rect 7969 35878 7983 35930
rect 7983 35878 7995 35930
rect 7995 35878 8025 35930
rect 8049 35878 8059 35930
rect 8059 35878 8105 35930
rect 7809 35876 7865 35878
rect 7889 35876 7945 35878
rect 7969 35876 8025 35878
rect 8049 35876 8105 35878
rect 7809 34842 7865 34844
rect 7889 34842 7945 34844
rect 7969 34842 8025 34844
rect 8049 34842 8105 34844
rect 7809 34790 7855 34842
rect 7855 34790 7865 34842
rect 7889 34790 7919 34842
rect 7919 34790 7931 34842
rect 7931 34790 7945 34842
rect 7969 34790 7983 34842
rect 7983 34790 7995 34842
rect 7995 34790 8025 34842
rect 8049 34790 8059 34842
rect 8059 34790 8105 34842
rect 7809 34788 7865 34790
rect 7889 34788 7945 34790
rect 7969 34788 8025 34790
rect 8049 34788 8105 34790
rect 7809 33754 7865 33756
rect 7889 33754 7945 33756
rect 7969 33754 8025 33756
rect 8049 33754 8105 33756
rect 7809 33702 7855 33754
rect 7855 33702 7865 33754
rect 7889 33702 7919 33754
rect 7919 33702 7931 33754
rect 7931 33702 7945 33754
rect 7969 33702 7983 33754
rect 7983 33702 7995 33754
rect 7995 33702 8025 33754
rect 8049 33702 8059 33754
rect 8059 33702 8105 33754
rect 7809 33700 7865 33702
rect 7889 33700 7945 33702
rect 7969 33700 8025 33702
rect 8049 33700 8105 33702
rect 7809 32666 7865 32668
rect 7889 32666 7945 32668
rect 7969 32666 8025 32668
rect 8049 32666 8105 32668
rect 7809 32614 7855 32666
rect 7855 32614 7865 32666
rect 7889 32614 7919 32666
rect 7919 32614 7931 32666
rect 7931 32614 7945 32666
rect 7969 32614 7983 32666
rect 7983 32614 7995 32666
rect 7995 32614 8025 32666
rect 8049 32614 8059 32666
rect 8059 32614 8105 32666
rect 7809 32612 7865 32614
rect 7889 32612 7945 32614
rect 7969 32612 8025 32614
rect 8049 32612 8105 32614
rect 7809 31578 7865 31580
rect 7889 31578 7945 31580
rect 7969 31578 8025 31580
rect 8049 31578 8105 31580
rect 7809 31526 7855 31578
rect 7855 31526 7865 31578
rect 7889 31526 7919 31578
rect 7919 31526 7931 31578
rect 7931 31526 7945 31578
rect 7969 31526 7983 31578
rect 7983 31526 7995 31578
rect 7995 31526 8025 31578
rect 8049 31526 8059 31578
rect 8059 31526 8105 31578
rect 7809 31524 7865 31526
rect 7889 31524 7945 31526
rect 7969 31524 8025 31526
rect 8049 31524 8105 31526
rect 7809 30490 7865 30492
rect 7889 30490 7945 30492
rect 7969 30490 8025 30492
rect 8049 30490 8105 30492
rect 7809 30438 7855 30490
rect 7855 30438 7865 30490
rect 7889 30438 7919 30490
rect 7919 30438 7931 30490
rect 7931 30438 7945 30490
rect 7969 30438 7983 30490
rect 7983 30438 7995 30490
rect 7995 30438 8025 30490
rect 8049 30438 8059 30490
rect 8059 30438 8105 30490
rect 7809 30436 7865 30438
rect 7889 30436 7945 30438
rect 7969 30436 8025 30438
rect 8049 30436 8105 30438
rect 7809 29402 7865 29404
rect 7889 29402 7945 29404
rect 7969 29402 8025 29404
rect 8049 29402 8105 29404
rect 7809 29350 7855 29402
rect 7855 29350 7865 29402
rect 7889 29350 7919 29402
rect 7919 29350 7931 29402
rect 7931 29350 7945 29402
rect 7969 29350 7983 29402
rect 7983 29350 7995 29402
rect 7995 29350 8025 29402
rect 8049 29350 8059 29402
rect 8059 29350 8105 29402
rect 7809 29348 7865 29350
rect 7889 29348 7945 29350
rect 7969 29348 8025 29350
rect 8049 29348 8105 29350
rect 8206 29280 8262 29336
rect 7809 28314 7865 28316
rect 7889 28314 7945 28316
rect 7969 28314 8025 28316
rect 8049 28314 8105 28316
rect 7809 28262 7855 28314
rect 7855 28262 7865 28314
rect 7889 28262 7919 28314
rect 7919 28262 7931 28314
rect 7931 28262 7945 28314
rect 7969 28262 7983 28314
rect 7983 28262 7995 28314
rect 7995 28262 8025 28314
rect 8049 28262 8059 28314
rect 8059 28262 8105 28314
rect 7809 28260 7865 28262
rect 7889 28260 7945 28262
rect 7969 28260 8025 28262
rect 8049 28260 8105 28262
rect 7809 27226 7865 27228
rect 7889 27226 7945 27228
rect 7969 27226 8025 27228
rect 8049 27226 8105 27228
rect 7809 27174 7855 27226
rect 7855 27174 7865 27226
rect 7889 27174 7919 27226
rect 7919 27174 7931 27226
rect 7931 27174 7945 27226
rect 7969 27174 7983 27226
rect 7983 27174 7995 27226
rect 7995 27174 8025 27226
rect 8049 27174 8059 27226
rect 8059 27174 8105 27226
rect 7809 27172 7865 27174
rect 7889 27172 7945 27174
rect 7969 27172 8025 27174
rect 8049 27172 8105 27174
rect 7809 26138 7865 26140
rect 7889 26138 7945 26140
rect 7969 26138 8025 26140
rect 8049 26138 8105 26140
rect 7809 26086 7855 26138
rect 7855 26086 7865 26138
rect 7889 26086 7919 26138
rect 7919 26086 7931 26138
rect 7931 26086 7945 26138
rect 7969 26086 7983 26138
rect 7983 26086 7995 26138
rect 7995 26086 8025 26138
rect 8049 26086 8059 26138
rect 8059 26086 8105 26138
rect 7809 26084 7865 26086
rect 7889 26084 7945 26086
rect 7969 26084 8025 26086
rect 8049 26084 8105 26086
rect 8206 25236 8208 25256
rect 8208 25236 8260 25256
rect 8260 25236 8262 25256
rect 8206 25200 8262 25236
rect 7809 25050 7865 25052
rect 7889 25050 7945 25052
rect 7969 25050 8025 25052
rect 8049 25050 8105 25052
rect 7809 24998 7855 25050
rect 7855 24998 7865 25050
rect 7889 24998 7919 25050
rect 7919 24998 7931 25050
rect 7931 24998 7945 25050
rect 7969 24998 7983 25050
rect 7983 24998 7995 25050
rect 7995 24998 8025 25050
rect 8049 24998 8059 25050
rect 8059 24998 8105 25050
rect 7809 24996 7865 24998
rect 7889 24996 7945 24998
rect 7969 24996 8025 24998
rect 8049 24996 8105 24998
rect 7010 20848 7066 20904
rect 6458 17604 6514 17640
rect 6458 17584 6460 17604
rect 6460 17584 6512 17604
rect 6512 17584 6514 17604
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 7562 21972 7564 21992
rect 7564 21972 7616 21992
rect 7616 21972 7618 21992
rect 7562 21936 7618 21972
rect 7378 18808 7434 18864
rect 7102 14320 7158 14376
rect 7102 13640 7158 13696
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 6826 10548 6828 10568
rect 6828 10548 6880 10568
rect 6880 10548 6882 10568
rect 6826 10512 6882 10548
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 7102 8916 7104 8936
rect 7104 8916 7156 8936
rect 7156 8916 7158 8936
rect 7102 8880 7158 8916
rect 7809 23962 7865 23964
rect 7889 23962 7945 23964
rect 7969 23962 8025 23964
rect 8049 23962 8105 23964
rect 7809 23910 7855 23962
rect 7855 23910 7865 23962
rect 7889 23910 7919 23962
rect 7919 23910 7931 23962
rect 7931 23910 7945 23962
rect 7969 23910 7983 23962
rect 7983 23910 7995 23962
rect 7995 23910 8025 23962
rect 8049 23910 8059 23962
rect 8059 23910 8105 23962
rect 7809 23908 7865 23910
rect 7889 23908 7945 23910
rect 7969 23908 8025 23910
rect 8049 23908 8105 23910
rect 7809 22874 7865 22876
rect 7889 22874 7945 22876
rect 7969 22874 8025 22876
rect 8049 22874 8105 22876
rect 7809 22822 7855 22874
rect 7855 22822 7865 22874
rect 7889 22822 7919 22874
rect 7919 22822 7931 22874
rect 7931 22822 7945 22874
rect 7969 22822 7983 22874
rect 7983 22822 7995 22874
rect 7995 22822 8025 22874
rect 8049 22822 8059 22874
rect 8059 22822 8105 22874
rect 7809 22820 7865 22822
rect 7889 22820 7945 22822
rect 7969 22820 8025 22822
rect 8049 22820 8105 22822
rect 7809 21786 7865 21788
rect 7889 21786 7945 21788
rect 7969 21786 8025 21788
rect 8049 21786 8105 21788
rect 7809 21734 7855 21786
rect 7855 21734 7865 21786
rect 7889 21734 7919 21786
rect 7919 21734 7931 21786
rect 7931 21734 7945 21786
rect 7969 21734 7983 21786
rect 7983 21734 7995 21786
rect 7995 21734 8025 21786
rect 8049 21734 8059 21786
rect 8059 21734 8105 21786
rect 7809 21732 7865 21734
rect 7889 21732 7945 21734
rect 7969 21732 8025 21734
rect 8049 21732 8105 21734
rect 9523 35386 9579 35388
rect 9603 35386 9659 35388
rect 9683 35386 9739 35388
rect 9763 35386 9819 35388
rect 9523 35334 9569 35386
rect 9569 35334 9579 35386
rect 9603 35334 9633 35386
rect 9633 35334 9645 35386
rect 9645 35334 9659 35386
rect 9683 35334 9697 35386
rect 9697 35334 9709 35386
rect 9709 35334 9739 35386
rect 9763 35334 9773 35386
rect 9773 35334 9819 35386
rect 9523 35332 9579 35334
rect 9603 35332 9659 35334
rect 9683 35332 9739 35334
rect 9763 35332 9819 35334
rect 9523 34298 9579 34300
rect 9603 34298 9659 34300
rect 9683 34298 9739 34300
rect 9763 34298 9819 34300
rect 9523 34246 9569 34298
rect 9569 34246 9579 34298
rect 9603 34246 9633 34298
rect 9633 34246 9645 34298
rect 9645 34246 9659 34298
rect 9683 34246 9697 34298
rect 9697 34246 9709 34298
rect 9709 34246 9739 34298
rect 9763 34246 9773 34298
rect 9773 34246 9819 34298
rect 9523 34244 9579 34246
rect 9603 34244 9659 34246
rect 9683 34244 9739 34246
rect 9763 34244 9819 34246
rect 10046 36216 10102 36272
rect 9523 33210 9579 33212
rect 9603 33210 9659 33212
rect 9683 33210 9739 33212
rect 9763 33210 9819 33212
rect 9523 33158 9569 33210
rect 9569 33158 9579 33210
rect 9603 33158 9633 33210
rect 9633 33158 9645 33210
rect 9645 33158 9659 33210
rect 9683 33158 9697 33210
rect 9697 33158 9709 33210
rect 9709 33158 9739 33210
rect 9763 33158 9773 33210
rect 9773 33158 9819 33210
rect 9523 33156 9579 33158
rect 9603 33156 9659 33158
rect 9683 33156 9739 33158
rect 9763 33156 9819 33158
rect 11236 37018 11292 37020
rect 11316 37018 11372 37020
rect 11396 37018 11452 37020
rect 11476 37018 11532 37020
rect 11236 36966 11282 37018
rect 11282 36966 11292 37018
rect 11316 36966 11346 37018
rect 11346 36966 11358 37018
rect 11358 36966 11372 37018
rect 11396 36966 11410 37018
rect 11410 36966 11422 37018
rect 11422 36966 11452 37018
rect 11476 36966 11486 37018
rect 11486 36966 11532 37018
rect 11236 36964 11292 36966
rect 11316 36964 11372 36966
rect 11396 36964 11452 36966
rect 11476 36964 11532 36966
rect 10506 35944 10562 36000
rect 10506 34992 10562 35048
rect 8574 29708 8630 29744
rect 8574 29688 8576 29708
rect 8576 29688 8628 29708
rect 8628 29688 8630 29708
rect 9523 32122 9579 32124
rect 9603 32122 9659 32124
rect 9683 32122 9739 32124
rect 9763 32122 9819 32124
rect 9523 32070 9569 32122
rect 9569 32070 9579 32122
rect 9603 32070 9633 32122
rect 9633 32070 9645 32122
rect 9645 32070 9659 32122
rect 9683 32070 9697 32122
rect 9697 32070 9709 32122
rect 9709 32070 9739 32122
rect 9763 32070 9773 32122
rect 9773 32070 9819 32122
rect 9523 32068 9579 32070
rect 9603 32068 9659 32070
rect 9683 32068 9739 32070
rect 9763 32068 9819 32070
rect 9523 31034 9579 31036
rect 9603 31034 9659 31036
rect 9683 31034 9739 31036
rect 9763 31034 9819 31036
rect 9523 30982 9569 31034
rect 9569 30982 9579 31034
rect 9603 30982 9633 31034
rect 9633 30982 9645 31034
rect 9645 30982 9659 31034
rect 9683 30982 9697 31034
rect 9697 30982 9709 31034
rect 9709 30982 9739 31034
rect 9763 30982 9773 31034
rect 9773 30982 9819 31034
rect 9523 30980 9579 30982
rect 9603 30980 9659 30982
rect 9683 30980 9739 30982
rect 9763 30980 9819 30982
rect 9218 29280 9274 29336
rect 8390 22636 8446 22672
rect 8390 22616 8392 22636
rect 8392 22616 8444 22636
rect 8444 22616 8446 22636
rect 7809 20698 7865 20700
rect 7889 20698 7945 20700
rect 7969 20698 8025 20700
rect 8049 20698 8105 20700
rect 7809 20646 7855 20698
rect 7855 20646 7865 20698
rect 7889 20646 7919 20698
rect 7919 20646 7931 20698
rect 7931 20646 7945 20698
rect 7969 20646 7983 20698
rect 7983 20646 7995 20698
rect 7995 20646 8025 20698
rect 8049 20646 8059 20698
rect 8059 20646 8105 20698
rect 7809 20644 7865 20646
rect 7889 20644 7945 20646
rect 7969 20644 8025 20646
rect 8049 20644 8105 20646
rect 7809 19610 7865 19612
rect 7889 19610 7945 19612
rect 7969 19610 8025 19612
rect 8049 19610 8105 19612
rect 7809 19558 7855 19610
rect 7855 19558 7865 19610
rect 7889 19558 7919 19610
rect 7919 19558 7931 19610
rect 7931 19558 7945 19610
rect 7969 19558 7983 19610
rect 7983 19558 7995 19610
rect 7995 19558 8025 19610
rect 8049 19558 8059 19610
rect 8059 19558 8105 19610
rect 7809 19556 7865 19558
rect 7889 19556 7945 19558
rect 7969 19556 8025 19558
rect 8049 19556 8105 19558
rect 7654 18672 7710 18728
rect 7838 18944 7894 19000
rect 7562 16496 7618 16552
rect 7809 18522 7865 18524
rect 7889 18522 7945 18524
rect 7969 18522 8025 18524
rect 8049 18522 8105 18524
rect 7809 18470 7855 18522
rect 7855 18470 7865 18522
rect 7889 18470 7919 18522
rect 7919 18470 7931 18522
rect 7931 18470 7945 18522
rect 7969 18470 7983 18522
rect 7983 18470 7995 18522
rect 7995 18470 8025 18522
rect 8049 18470 8059 18522
rect 8059 18470 8105 18522
rect 7809 18468 7865 18470
rect 7889 18468 7945 18470
rect 7969 18468 8025 18470
rect 8049 18468 8105 18470
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 8666 24268 8722 24304
rect 8666 24248 8668 24268
rect 8668 24248 8720 24268
rect 8720 24248 8722 24268
rect 8850 23060 8852 23080
rect 8852 23060 8904 23080
rect 8904 23060 8906 23080
rect 8850 23024 8906 23060
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 8206 15156 8262 15192
rect 8206 15136 8208 15156
rect 8208 15136 8260 15156
rect 8260 15136 8262 15156
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 7470 11636 7472 11656
rect 7472 11636 7524 11656
rect 7524 11636 7526 11656
rect 7470 11600 7526 11636
rect 8114 12824 8170 12880
rect 7746 12144 7802 12200
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 7194 8472 7250 8528
rect 2669 1658 2725 1660
rect 2749 1658 2805 1660
rect 2829 1658 2885 1660
rect 2909 1658 2965 1660
rect 2669 1606 2715 1658
rect 2715 1606 2725 1658
rect 2749 1606 2779 1658
rect 2779 1606 2791 1658
rect 2791 1606 2805 1658
rect 2829 1606 2843 1658
rect 2843 1606 2855 1658
rect 2855 1606 2885 1658
rect 2909 1606 2919 1658
rect 2919 1606 2965 1658
rect 2669 1604 2725 1606
rect 2749 1604 2805 1606
rect 2829 1604 2885 1606
rect 2909 1604 2965 1606
rect 6096 1658 6152 1660
rect 6176 1658 6232 1660
rect 6256 1658 6312 1660
rect 6336 1658 6392 1660
rect 6096 1606 6142 1658
rect 6142 1606 6152 1658
rect 6176 1606 6206 1658
rect 6206 1606 6218 1658
rect 6218 1606 6232 1658
rect 6256 1606 6270 1658
rect 6270 1606 6282 1658
rect 6282 1606 6312 1658
rect 6336 1606 6346 1658
rect 6346 1606 6392 1658
rect 6096 1604 6152 1606
rect 6176 1604 6232 1606
rect 6256 1604 6312 1606
rect 6336 1604 6392 1606
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 8482 10512 8538 10568
rect 8298 5752 8354 5808
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 9218 28464 9274 28520
rect 9523 29946 9579 29948
rect 9603 29946 9659 29948
rect 9683 29946 9739 29948
rect 9763 29946 9819 29948
rect 9523 29894 9569 29946
rect 9569 29894 9579 29946
rect 9603 29894 9633 29946
rect 9633 29894 9645 29946
rect 9645 29894 9659 29946
rect 9683 29894 9697 29946
rect 9697 29894 9709 29946
rect 9709 29894 9739 29946
rect 9763 29894 9773 29946
rect 9773 29894 9819 29946
rect 9523 29892 9579 29894
rect 9603 29892 9659 29894
rect 9683 29892 9739 29894
rect 9763 29892 9819 29894
rect 9586 29688 9642 29744
rect 10690 34584 10746 34640
rect 10966 36080 11022 36136
rect 11236 35930 11292 35932
rect 11316 35930 11372 35932
rect 11396 35930 11452 35932
rect 11476 35930 11532 35932
rect 11236 35878 11282 35930
rect 11282 35878 11292 35930
rect 11316 35878 11346 35930
rect 11346 35878 11358 35930
rect 11358 35878 11372 35930
rect 11396 35878 11410 35930
rect 11410 35878 11422 35930
rect 11422 35878 11452 35930
rect 11476 35878 11486 35930
rect 11486 35878 11532 35930
rect 11236 35876 11292 35878
rect 11316 35876 11372 35878
rect 11396 35876 11452 35878
rect 11476 35876 11532 35878
rect 9523 28858 9579 28860
rect 9603 28858 9659 28860
rect 9683 28858 9739 28860
rect 9763 28858 9819 28860
rect 9523 28806 9569 28858
rect 9569 28806 9579 28858
rect 9603 28806 9633 28858
rect 9633 28806 9645 28858
rect 9645 28806 9659 28858
rect 9683 28806 9697 28858
rect 9697 28806 9709 28858
rect 9709 28806 9739 28858
rect 9763 28806 9773 28858
rect 9773 28806 9819 28858
rect 9523 28804 9579 28806
rect 9603 28804 9659 28806
rect 9683 28804 9739 28806
rect 9763 28804 9819 28806
rect 9586 28056 9642 28112
rect 9523 27770 9579 27772
rect 9603 27770 9659 27772
rect 9683 27770 9739 27772
rect 9763 27770 9819 27772
rect 9523 27718 9569 27770
rect 9569 27718 9579 27770
rect 9603 27718 9633 27770
rect 9633 27718 9645 27770
rect 9645 27718 9659 27770
rect 9683 27718 9697 27770
rect 9697 27718 9709 27770
rect 9709 27718 9739 27770
rect 9763 27718 9773 27770
rect 9773 27718 9819 27770
rect 9523 27716 9579 27718
rect 9603 27716 9659 27718
rect 9683 27716 9739 27718
rect 9763 27716 9819 27718
rect 9862 27376 9918 27432
rect 9523 26682 9579 26684
rect 9603 26682 9659 26684
rect 9683 26682 9739 26684
rect 9763 26682 9819 26684
rect 9523 26630 9569 26682
rect 9569 26630 9579 26682
rect 9603 26630 9633 26682
rect 9633 26630 9645 26682
rect 9645 26630 9659 26682
rect 9683 26630 9697 26682
rect 9697 26630 9709 26682
rect 9709 26630 9739 26682
rect 9763 26630 9773 26682
rect 9773 26630 9819 26682
rect 9523 26628 9579 26630
rect 9603 26628 9659 26630
rect 9683 26628 9739 26630
rect 9763 26628 9819 26630
rect 9523 25594 9579 25596
rect 9603 25594 9659 25596
rect 9683 25594 9739 25596
rect 9763 25594 9819 25596
rect 9523 25542 9569 25594
rect 9569 25542 9579 25594
rect 9603 25542 9633 25594
rect 9633 25542 9645 25594
rect 9645 25542 9659 25594
rect 9683 25542 9697 25594
rect 9697 25542 9709 25594
rect 9709 25542 9739 25594
rect 9763 25542 9773 25594
rect 9773 25542 9819 25594
rect 9523 25540 9579 25542
rect 9603 25540 9659 25542
rect 9683 25540 9739 25542
rect 9763 25540 9819 25542
rect 9523 24506 9579 24508
rect 9603 24506 9659 24508
rect 9683 24506 9739 24508
rect 9763 24506 9819 24508
rect 9523 24454 9569 24506
rect 9569 24454 9579 24506
rect 9603 24454 9633 24506
rect 9633 24454 9645 24506
rect 9645 24454 9659 24506
rect 9683 24454 9697 24506
rect 9697 24454 9709 24506
rect 9709 24454 9739 24506
rect 9763 24454 9773 24506
rect 9773 24454 9819 24506
rect 9523 24452 9579 24454
rect 9603 24452 9659 24454
rect 9683 24452 9739 24454
rect 9763 24452 9819 24454
rect 9494 24248 9550 24304
rect 8942 20848 8998 20904
rect 9523 23418 9579 23420
rect 9603 23418 9659 23420
rect 9683 23418 9739 23420
rect 9763 23418 9819 23420
rect 9523 23366 9569 23418
rect 9569 23366 9579 23418
rect 9603 23366 9633 23418
rect 9633 23366 9645 23418
rect 9645 23366 9659 23418
rect 9683 23366 9697 23418
rect 9697 23366 9709 23418
rect 9709 23366 9739 23418
rect 9763 23366 9773 23418
rect 9773 23366 9819 23418
rect 9523 23364 9579 23366
rect 9603 23364 9659 23366
rect 9683 23364 9739 23366
rect 9763 23364 9819 23366
rect 9523 22330 9579 22332
rect 9603 22330 9659 22332
rect 9683 22330 9739 22332
rect 9763 22330 9819 22332
rect 9523 22278 9569 22330
rect 9569 22278 9579 22330
rect 9603 22278 9633 22330
rect 9633 22278 9645 22330
rect 9645 22278 9659 22330
rect 9683 22278 9697 22330
rect 9697 22278 9709 22330
rect 9709 22278 9739 22330
rect 9763 22278 9773 22330
rect 9773 22278 9819 22330
rect 9523 22276 9579 22278
rect 9603 22276 9659 22278
rect 9683 22276 9739 22278
rect 9763 22276 9819 22278
rect 9862 21936 9918 21992
rect 9770 21664 9826 21720
rect 10138 26288 10194 26344
rect 9523 21242 9579 21244
rect 9603 21242 9659 21244
rect 9683 21242 9739 21244
rect 9763 21242 9819 21244
rect 9523 21190 9569 21242
rect 9569 21190 9579 21242
rect 9603 21190 9633 21242
rect 9633 21190 9645 21242
rect 9645 21190 9659 21242
rect 9683 21190 9697 21242
rect 9697 21190 9709 21242
rect 9709 21190 9739 21242
rect 9763 21190 9773 21242
rect 9773 21190 9819 21242
rect 9523 21188 9579 21190
rect 9603 21188 9659 21190
rect 9683 21188 9739 21190
rect 9763 21188 9819 21190
rect 9034 19508 9090 19544
rect 9034 19488 9036 19508
rect 9036 19488 9088 19508
rect 9088 19488 9090 19508
rect 8942 16108 8998 16144
rect 8942 16088 8944 16108
rect 8944 16088 8996 16108
rect 8996 16088 8998 16108
rect 9523 20154 9579 20156
rect 9603 20154 9659 20156
rect 9683 20154 9739 20156
rect 9763 20154 9819 20156
rect 9523 20102 9569 20154
rect 9569 20102 9579 20154
rect 9603 20102 9633 20154
rect 9633 20102 9645 20154
rect 9645 20102 9659 20154
rect 9683 20102 9697 20154
rect 9697 20102 9709 20154
rect 9709 20102 9739 20154
rect 9763 20102 9773 20154
rect 9773 20102 9819 20154
rect 9523 20100 9579 20102
rect 9603 20100 9659 20102
rect 9683 20100 9739 20102
rect 9763 20100 9819 20102
rect 9954 20032 10010 20088
rect 10138 20032 10194 20088
rect 11236 34842 11292 34844
rect 11316 34842 11372 34844
rect 11396 34842 11452 34844
rect 11476 34842 11532 34844
rect 11236 34790 11282 34842
rect 11282 34790 11292 34842
rect 11316 34790 11346 34842
rect 11346 34790 11358 34842
rect 11358 34790 11372 34842
rect 11396 34790 11410 34842
rect 11410 34790 11422 34842
rect 11422 34790 11452 34842
rect 11476 34790 11486 34842
rect 11486 34790 11532 34842
rect 11236 34788 11292 34790
rect 11316 34788 11372 34790
rect 11396 34788 11452 34790
rect 11476 34788 11532 34790
rect 11518 33940 11520 33960
rect 11520 33940 11572 33960
rect 11572 33940 11574 33960
rect 11518 33904 11574 33940
rect 12950 38650 13006 38652
rect 13030 38650 13086 38652
rect 13110 38650 13166 38652
rect 13190 38650 13246 38652
rect 12950 38598 12996 38650
rect 12996 38598 13006 38650
rect 13030 38598 13060 38650
rect 13060 38598 13072 38650
rect 13072 38598 13086 38650
rect 13110 38598 13124 38650
rect 13124 38598 13136 38650
rect 13136 38598 13166 38650
rect 13190 38598 13200 38650
rect 13200 38598 13246 38650
rect 12950 38596 13006 38598
rect 13030 38596 13086 38598
rect 13110 38596 13166 38598
rect 13190 38596 13246 38598
rect 13910 38936 13966 38992
rect 13634 38392 13690 38448
rect 12950 37562 13006 37564
rect 13030 37562 13086 37564
rect 13110 37562 13166 37564
rect 13190 37562 13246 37564
rect 12950 37510 12996 37562
rect 12996 37510 13006 37562
rect 13030 37510 13060 37562
rect 13060 37510 13072 37562
rect 13072 37510 13086 37562
rect 13110 37510 13124 37562
rect 13124 37510 13136 37562
rect 13136 37510 13166 37562
rect 13190 37510 13200 37562
rect 13200 37510 13246 37562
rect 12950 37508 13006 37510
rect 13030 37508 13086 37510
rect 13110 37508 13166 37510
rect 13190 37508 13246 37510
rect 13082 37204 13084 37224
rect 13084 37204 13136 37224
rect 13136 37204 13138 37224
rect 13082 37168 13138 37204
rect 12950 36474 13006 36476
rect 13030 36474 13086 36476
rect 13110 36474 13166 36476
rect 13190 36474 13246 36476
rect 12950 36422 12996 36474
rect 12996 36422 13006 36474
rect 13030 36422 13060 36474
rect 13060 36422 13072 36474
rect 13072 36422 13086 36474
rect 13110 36422 13124 36474
rect 13124 36422 13136 36474
rect 13136 36422 13166 36474
rect 13190 36422 13200 36474
rect 13200 36422 13246 36474
rect 12950 36420 13006 36422
rect 13030 36420 13086 36422
rect 13110 36420 13166 36422
rect 13190 36420 13246 36422
rect 14186 38528 14242 38584
rect 13818 37848 13874 37904
rect 13450 36624 13506 36680
rect 14002 37304 14058 37360
rect 12530 35128 12586 35184
rect 11236 33754 11292 33756
rect 11316 33754 11372 33756
rect 11396 33754 11452 33756
rect 11476 33754 11532 33756
rect 11236 33702 11282 33754
rect 11282 33702 11292 33754
rect 11316 33702 11346 33754
rect 11346 33702 11358 33754
rect 11358 33702 11372 33754
rect 11396 33702 11410 33754
rect 11410 33702 11422 33754
rect 11422 33702 11452 33754
rect 11476 33702 11486 33754
rect 11486 33702 11532 33754
rect 11236 33700 11292 33702
rect 11316 33700 11372 33702
rect 11396 33700 11452 33702
rect 11476 33700 11532 33702
rect 11058 31864 11114 31920
rect 10782 29960 10838 30016
rect 10690 29844 10746 29880
rect 10690 29824 10692 29844
rect 10692 29824 10744 29844
rect 10744 29824 10746 29844
rect 10414 25064 10470 25120
rect 9862 19624 9918 19680
rect 10138 19624 10194 19680
rect 9523 19066 9579 19068
rect 9603 19066 9659 19068
rect 9683 19066 9739 19068
rect 9763 19066 9819 19068
rect 9523 19014 9569 19066
rect 9569 19014 9579 19066
rect 9603 19014 9633 19066
rect 9633 19014 9645 19066
rect 9645 19014 9659 19066
rect 9683 19014 9697 19066
rect 9697 19014 9709 19066
rect 9709 19014 9739 19066
rect 9763 19014 9773 19066
rect 9773 19014 9819 19066
rect 9523 19012 9579 19014
rect 9603 19012 9659 19014
rect 9683 19012 9739 19014
rect 9763 19012 9819 19014
rect 9586 18808 9642 18864
rect 10046 19488 10102 19544
rect 9678 18672 9734 18728
rect 9523 17978 9579 17980
rect 9603 17978 9659 17980
rect 9683 17978 9739 17980
rect 9763 17978 9819 17980
rect 9523 17926 9569 17978
rect 9569 17926 9579 17978
rect 9603 17926 9633 17978
rect 9633 17926 9645 17978
rect 9645 17926 9659 17978
rect 9683 17926 9697 17978
rect 9697 17926 9709 17978
rect 9709 17926 9739 17978
rect 9763 17926 9773 17978
rect 9773 17926 9819 17978
rect 9523 17924 9579 17926
rect 9603 17924 9659 17926
rect 9683 17924 9739 17926
rect 9763 17924 9819 17926
rect 9678 17720 9734 17776
rect 9678 17040 9734 17096
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 9218 16496 9274 16552
rect 8850 11600 8906 11656
rect 9310 16088 9366 16144
rect 9034 13948 9036 13968
rect 9036 13948 9088 13968
rect 9088 13948 9090 13968
rect 9034 13912 9090 13948
rect 10138 17992 10194 18048
rect 9954 16360 10010 16416
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 10138 16768 10194 16824
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 8850 10648 8906 10704
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 9034 6704 9090 6760
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 9954 13912 10010 13968
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 11236 32666 11292 32668
rect 11316 32666 11372 32668
rect 11396 32666 11452 32668
rect 11476 32666 11532 32668
rect 11236 32614 11282 32666
rect 11282 32614 11292 32666
rect 11316 32614 11346 32666
rect 11346 32614 11358 32666
rect 11358 32614 11372 32666
rect 11396 32614 11410 32666
rect 11410 32614 11422 32666
rect 11422 32614 11452 32666
rect 11476 32614 11486 32666
rect 11486 32614 11532 32666
rect 11236 32612 11292 32614
rect 11316 32612 11372 32614
rect 11396 32612 11452 32614
rect 11476 32612 11532 32614
rect 11518 31864 11574 31920
rect 11236 31578 11292 31580
rect 11316 31578 11372 31580
rect 11396 31578 11452 31580
rect 11476 31578 11532 31580
rect 11236 31526 11282 31578
rect 11282 31526 11292 31578
rect 11316 31526 11346 31578
rect 11346 31526 11358 31578
rect 11358 31526 11372 31578
rect 11396 31526 11410 31578
rect 11410 31526 11422 31578
rect 11422 31526 11452 31578
rect 11476 31526 11486 31578
rect 11486 31526 11532 31578
rect 11236 31524 11292 31526
rect 11316 31524 11372 31526
rect 11396 31524 11452 31526
rect 11476 31524 11532 31526
rect 11242 30776 11298 30832
rect 11236 30490 11292 30492
rect 11316 30490 11372 30492
rect 11396 30490 11452 30492
rect 11476 30490 11532 30492
rect 11236 30438 11282 30490
rect 11282 30438 11292 30490
rect 11316 30438 11346 30490
rect 11346 30438 11358 30490
rect 11358 30438 11372 30490
rect 11396 30438 11410 30490
rect 11410 30438 11422 30490
rect 11422 30438 11452 30490
rect 11476 30438 11486 30490
rect 11486 30438 11532 30490
rect 11236 30436 11292 30438
rect 11316 30436 11372 30438
rect 11396 30436 11452 30438
rect 11476 30436 11532 30438
rect 11150 29960 11206 30016
rect 11610 30232 11666 30288
rect 11058 28736 11114 28792
rect 11058 28464 11114 28520
rect 11334 29960 11390 30016
rect 11426 29824 11482 29880
rect 11242 29688 11298 29744
rect 11242 29588 11244 29608
rect 11244 29588 11296 29608
rect 11296 29588 11298 29608
rect 11242 29552 11298 29588
rect 11236 29402 11292 29404
rect 11316 29402 11372 29404
rect 11396 29402 11452 29404
rect 11476 29402 11532 29404
rect 11236 29350 11282 29402
rect 11282 29350 11292 29402
rect 11316 29350 11346 29402
rect 11346 29350 11358 29402
rect 11358 29350 11372 29402
rect 11396 29350 11410 29402
rect 11410 29350 11422 29402
rect 11422 29350 11452 29402
rect 11476 29350 11486 29402
rect 11486 29350 11532 29402
rect 11236 29348 11292 29350
rect 11316 29348 11372 29350
rect 11396 29348 11452 29350
rect 11476 29348 11532 29350
rect 11610 29008 11666 29064
rect 11236 28314 11292 28316
rect 11316 28314 11372 28316
rect 11396 28314 11452 28316
rect 11476 28314 11532 28316
rect 11236 28262 11282 28314
rect 11282 28262 11292 28314
rect 11316 28262 11346 28314
rect 11346 28262 11358 28314
rect 11358 28262 11372 28314
rect 11396 28262 11410 28314
rect 11410 28262 11422 28314
rect 11422 28262 11452 28314
rect 11476 28262 11486 28314
rect 11486 28262 11532 28314
rect 11236 28260 11292 28262
rect 11316 28260 11372 28262
rect 11396 28260 11452 28262
rect 11476 28260 11532 28262
rect 10414 17856 10470 17912
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 9862 8492 9918 8528
rect 9862 8472 9864 8492
rect 9864 8472 9916 8492
rect 9916 8472 9918 8492
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 10322 10512 10378 10568
rect 10138 8916 10140 8936
rect 10140 8916 10192 8936
rect 10192 8916 10194 8936
rect 10138 8880 10194 8916
rect 9678 6196 9680 6216
rect 9680 6196 9732 6216
rect 9732 6196 9734 6216
rect 9678 6160 9734 6196
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 11518 27376 11574 27432
rect 11236 27226 11292 27228
rect 11316 27226 11372 27228
rect 11396 27226 11452 27228
rect 11476 27226 11532 27228
rect 11236 27174 11282 27226
rect 11282 27174 11292 27226
rect 11316 27174 11346 27226
rect 11346 27174 11358 27226
rect 11358 27174 11372 27226
rect 11396 27174 11410 27226
rect 11410 27174 11422 27226
rect 11422 27174 11452 27226
rect 11476 27174 11486 27226
rect 11486 27174 11532 27226
rect 11236 27172 11292 27174
rect 11316 27172 11372 27174
rect 11396 27172 11452 27174
rect 11476 27172 11532 27174
rect 11236 26138 11292 26140
rect 11316 26138 11372 26140
rect 11396 26138 11452 26140
rect 11476 26138 11532 26140
rect 11236 26086 11282 26138
rect 11282 26086 11292 26138
rect 11316 26086 11346 26138
rect 11346 26086 11358 26138
rect 11358 26086 11372 26138
rect 11396 26086 11410 26138
rect 11410 26086 11422 26138
rect 11422 26086 11452 26138
rect 11476 26086 11486 26138
rect 11486 26086 11532 26138
rect 11236 26084 11292 26086
rect 11316 26084 11372 26086
rect 11396 26084 11452 26086
rect 11476 26084 11532 26086
rect 11150 25200 11206 25256
rect 11236 25050 11292 25052
rect 11316 25050 11372 25052
rect 11396 25050 11452 25052
rect 11476 25050 11532 25052
rect 11236 24998 11282 25050
rect 11282 24998 11292 25050
rect 11316 24998 11346 25050
rect 11346 24998 11358 25050
rect 11358 24998 11372 25050
rect 11396 24998 11410 25050
rect 11410 24998 11422 25050
rect 11422 24998 11452 25050
rect 11476 24998 11486 25050
rect 11486 24998 11532 25050
rect 11236 24996 11292 24998
rect 11316 24996 11372 24998
rect 11396 24996 11452 24998
rect 11476 24996 11532 24998
rect 12254 34448 12310 34504
rect 11978 31764 11980 31784
rect 11980 31764 12032 31784
rect 12032 31764 12034 31784
rect 11978 31728 12034 31764
rect 11886 31340 11942 31376
rect 11886 31320 11888 31340
rect 11888 31320 11940 31340
rect 11940 31320 11942 31340
rect 12162 33360 12218 33416
rect 12346 32408 12402 32464
rect 13266 36216 13322 36272
rect 13266 35672 13322 35728
rect 12950 35386 13006 35388
rect 13030 35386 13086 35388
rect 13110 35386 13166 35388
rect 13190 35386 13246 35388
rect 12950 35334 12996 35386
rect 12996 35334 13006 35386
rect 13030 35334 13060 35386
rect 13060 35334 13072 35386
rect 13072 35334 13086 35386
rect 13110 35334 13124 35386
rect 13124 35334 13136 35386
rect 13136 35334 13166 35386
rect 13190 35334 13200 35386
rect 13200 35334 13246 35386
rect 12950 35332 13006 35334
rect 13030 35332 13086 35334
rect 13110 35332 13166 35334
rect 13190 35332 13246 35334
rect 12950 34298 13006 34300
rect 13030 34298 13086 34300
rect 13110 34298 13166 34300
rect 13190 34298 13246 34300
rect 12950 34246 12996 34298
rect 12996 34246 13006 34298
rect 13030 34246 13060 34298
rect 13060 34246 13072 34298
rect 13072 34246 13086 34298
rect 13110 34246 13124 34298
rect 13124 34246 13136 34298
rect 13136 34246 13166 34298
rect 13190 34246 13200 34298
rect 13200 34246 13246 34298
rect 12950 34244 13006 34246
rect 13030 34244 13086 34246
rect 13110 34244 13166 34246
rect 13190 34244 13246 34246
rect 13266 34040 13322 34096
rect 12622 32544 12678 32600
rect 11794 29688 11850 29744
rect 12162 30776 12218 30832
rect 12346 31320 12402 31376
rect 12950 33210 13006 33212
rect 13030 33210 13086 33212
rect 13110 33210 13166 33212
rect 13190 33210 13246 33212
rect 12950 33158 12996 33210
rect 12996 33158 13006 33210
rect 13030 33158 13060 33210
rect 13060 33158 13072 33210
rect 13072 33158 13086 33210
rect 13110 33158 13124 33210
rect 13124 33158 13136 33210
rect 13136 33158 13166 33210
rect 13190 33158 13200 33210
rect 13200 33158 13246 33210
rect 12950 33156 13006 33158
rect 13030 33156 13086 33158
rect 13110 33156 13166 33158
rect 13190 33156 13246 33158
rect 12990 32272 13046 32328
rect 12950 32122 13006 32124
rect 13030 32122 13086 32124
rect 13110 32122 13166 32124
rect 13190 32122 13246 32124
rect 12950 32070 12996 32122
rect 12996 32070 13006 32122
rect 13030 32070 13060 32122
rect 13060 32070 13072 32122
rect 13072 32070 13086 32122
rect 13110 32070 13124 32122
rect 13124 32070 13136 32122
rect 13136 32070 13166 32122
rect 13190 32070 13200 32122
rect 13200 32070 13246 32122
rect 12950 32068 13006 32070
rect 13030 32068 13086 32070
rect 13110 32068 13166 32070
rect 13190 32068 13246 32070
rect 13726 36760 13782 36816
rect 13818 36216 13874 36272
rect 13726 36080 13782 36136
rect 13634 34992 13690 35048
rect 13542 34604 13598 34640
rect 13542 34584 13544 34604
rect 13544 34584 13596 34604
rect 13596 34584 13598 34604
rect 13358 33088 13414 33144
rect 13634 33632 13690 33688
rect 13818 34584 13874 34640
rect 14663 41370 14719 41372
rect 14743 41370 14799 41372
rect 14823 41370 14879 41372
rect 14903 41370 14959 41372
rect 14663 41318 14709 41370
rect 14709 41318 14719 41370
rect 14743 41318 14773 41370
rect 14773 41318 14785 41370
rect 14785 41318 14799 41370
rect 14823 41318 14837 41370
rect 14837 41318 14849 41370
rect 14849 41318 14879 41370
rect 14903 41318 14913 41370
rect 14913 41318 14959 41370
rect 14663 41316 14719 41318
rect 14743 41316 14799 41318
rect 14823 41316 14879 41318
rect 14903 41316 14959 41318
rect 14663 40282 14719 40284
rect 14743 40282 14799 40284
rect 14823 40282 14879 40284
rect 14903 40282 14959 40284
rect 14663 40230 14709 40282
rect 14709 40230 14719 40282
rect 14743 40230 14773 40282
rect 14773 40230 14785 40282
rect 14785 40230 14799 40282
rect 14823 40230 14837 40282
rect 14837 40230 14849 40282
rect 14849 40230 14879 40282
rect 14903 40230 14913 40282
rect 14913 40230 14959 40282
rect 14663 40228 14719 40230
rect 14743 40228 14799 40230
rect 14823 40228 14879 40230
rect 14903 40228 14959 40230
rect 14663 39194 14719 39196
rect 14743 39194 14799 39196
rect 14823 39194 14879 39196
rect 14903 39194 14959 39196
rect 14663 39142 14709 39194
rect 14709 39142 14719 39194
rect 14743 39142 14773 39194
rect 14773 39142 14785 39194
rect 14785 39142 14799 39194
rect 14823 39142 14837 39194
rect 14837 39142 14849 39194
rect 14849 39142 14879 39194
rect 14903 39142 14913 39194
rect 14913 39142 14959 39194
rect 14663 39140 14719 39142
rect 14743 39140 14799 39142
rect 14823 39140 14879 39142
rect 14903 39140 14959 39142
rect 14370 38664 14426 38720
rect 14663 38106 14719 38108
rect 14743 38106 14799 38108
rect 14823 38106 14879 38108
rect 14903 38106 14959 38108
rect 14663 38054 14709 38106
rect 14709 38054 14719 38106
rect 14743 38054 14773 38106
rect 14773 38054 14785 38106
rect 14785 38054 14799 38106
rect 14823 38054 14837 38106
rect 14837 38054 14849 38106
rect 14849 38054 14879 38106
rect 14903 38054 14913 38106
rect 14913 38054 14959 38106
rect 14663 38052 14719 38054
rect 14743 38052 14799 38054
rect 14823 38052 14879 38054
rect 14903 38052 14959 38054
rect 14370 37576 14426 37632
rect 14663 37018 14719 37020
rect 14743 37018 14799 37020
rect 14823 37018 14879 37020
rect 14903 37018 14959 37020
rect 14663 36966 14709 37018
rect 14709 36966 14719 37018
rect 14743 36966 14773 37018
rect 14773 36966 14785 37018
rect 14785 36966 14799 37018
rect 14823 36966 14837 37018
rect 14837 36966 14849 37018
rect 14849 36966 14879 37018
rect 14903 36966 14913 37018
rect 14913 36966 14959 37018
rect 14663 36964 14719 36966
rect 14743 36964 14799 36966
rect 14823 36964 14879 36966
rect 14903 36964 14959 36966
rect 14370 36488 14426 36544
rect 14663 35930 14719 35932
rect 14743 35930 14799 35932
rect 14823 35930 14879 35932
rect 14903 35930 14959 35932
rect 14663 35878 14709 35930
rect 14709 35878 14719 35930
rect 14743 35878 14773 35930
rect 14773 35878 14785 35930
rect 14785 35878 14799 35930
rect 14823 35878 14837 35930
rect 14837 35878 14849 35930
rect 14849 35878 14879 35930
rect 14903 35878 14913 35930
rect 14913 35878 14959 35930
rect 14663 35876 14719 35878
rect 14743 35876 14799 35878
rect 14823 35876 14879 35878
rect 14903 35876 14959 35878
rect 14462 35128 14518 35184
rect 13818 33224 13874 33280
rect 13634 32952 13690 33008
rect 13358 31184 13414 31240
rect 12950 31034 13006 31036
rect 13030 31034 13086 31036
rect 13110 31034 13166 31036
rect 13190 31034 13246 31036
rect 12950 30982 12996 31034
rect 12996 30982 13006 31034
rect 13030 30982 13060 31034
rect 13060 30982 13072 31034
rect 13072 30982 13086 31034
rect 13110 30982 13124 31034
rect 13124 30982 13136 31034
rect 13136 30982 13166 31034
rect 13190 30982 13200 31034
rect 13200 30982 13246 31034
rect 12950 30980 13006 30982
rect 13030 30980 13086 30982
rect 13110 30980 13166 30982
rect 13190 30980 13246 30982
rect 11236 23962 11292 23964
rect 11316 23962 11372 23964
rect 11396 23962 11452 23964
rect 11476 23962 11532 23964
rect 11236 23910 11282 23962
rect 11282 23910 11292 23962
rect 11316 23910 11346 23962
rect 11346 23910 11358 23962
rect 11358 23910 11372 23962
rect 11396 23910 11410 23962
rect 11410 23910 11422 23962
rect 11422 23910 11452 23962
rect 11476 23910 11486 23962
rect 11486 23910 11532 23962
rect 11236 23908 11292 23910
rect 11316 23908 11372 23910
rect 11396 23908 11452 23910
rect 11476 23908 11532 23910
rect 11236 22874 11292 22876
rect 11316 22874 11372 22876
rect 11396 22874 11452 22876
rect 11476 22874 11532 22876
rect 11236 22822 11282 22874
rect 11282 22822 11292 22874
rect 11316 22822 11346 22874
rect 11346 22822 11358 22874
rect 11358 22822 11372 22874
rect 11396 22822 11410 22874
rect 11410 22822 11422 22874
rect 11422 22822 11452 22874
rect 11476 22822 11486 22874
rect 11486 22822 11532 22874
rect 11236 22820 11292 22822
rect 11316 22820 11372 22822
rect 11396 22820 11452 22822
rect 11476 22820 11532 22822
rect 11150 22616 11206 22672
rect 12254 30096 12310 30152
rect 12346 29824 12402 29880
rect 12254 29144 12310 29200
rect 11978 27512 12034 27568
rect 12346 28056 12402 28112
rect 12622 29552 12678 29608
rect 12622 29008 12678 29064
rect 12950 29946 13006 29948
rect 13030 29946 13086 29948
rect 13110 29946 13166 29948
rect 13190 29946 13246 29948
rect 12950 29894 12996 29946
rect 12996 29894 13006 29946
rect 13030 29894 13060 29946
rect 13060 29894 13072 29946
rect 13072 29894 13086 29946
rect 13110 29894 13124 29946
rect 13124 29894 13136 29946
rect 13136 29894 13166 29946
rect 13190 29894 13200 29946
rect 13200 29894 13246 29946
rect 12950 29892 13006 29894
rect 13030 29892 13086 29894
rect 13110 29892 13166 29894
rect 13190 29892 13246 29894
rect 13174 29044 13176 29064
rect 13176 29044 13228 29064
rect 13228 29044 13230 29064
rect 13174 29008 13230 29044
rect 12950 28858 13006 28860
rect 13030 28858 13086 28860
rect 13110 28858 13166 28860
rect 13190 28858 13246 28860
rect 12950 28806 12996 28858
rect 12996 28806 13006 28858
rect 13030 28806 13060 28858
rect 13060 28806 13072 28858
rect 13072 28806 13086 28858
rect 13110 28806 13124 28858
rect 13124 28806 13136 28858
rect 13136 28806 13166 28858
rect 13190 28806 13200 28858
rect 13200 28806 13246 28858
rect 12950 28804 13006 28806
rect 13030 28804 13086 28806
rect 13110 28804 13166 28806
rect 13190 28804 13246 28806
rect 11886 26424 11942 26480
rect 11886 24792 11942 24848
rect 12254 25744 12310 25800
rect 11978 24248 12034 24304
rect 11236 21786 11292 21788
rect 11316 21786 11372 21788
rect 11396 21786 11452 21788
rect 11476 21786 11532 21788
rect 11236 21734 11282 21786
rect 11282 21734 11292 21786
rect 11316 21734 11346 21786
rect 11346 21734 11358 21786
rect 11358 21734 11372 21786
rect 11396 21734 11410 21786
rect 11410 21734 11422 21786
rect 11422 21734 11452 21786
rect 11476 21734 11486 21786
rect 11486 21734 11532 21786
rect 11236 21732 11292 21734
rect 11316 21732 11372 21734
rect 11396 21732 11452 21734
rect 11476 21732 11532 21734
rect 11236 20698 11292 20700
rect 11316 20698 11372 20700
rect 11396 20698 11452 20700
rect 11476 20698 11532 20700
rect 11236 20646 11282 20698
rect 11282 20646 11292 20698
rect 11316 20646 11346 20698
rect 11346 20646 11358 20698
rect 11358 20646 11372 20698
rect 11396 20646 11410 20698
rect 11410 20646 11422 20698
rect 11422 20646 11452 20698
rect 11476 20646 11486 20698
rect 11486 20646 11532 20698
rect 11236 20644 11292 20646
rect 11316 20644 11372 20646
rect 11396 20644 11452 20646
rect 11476 20644 11532 20646
rect 11794 21392 11850 21448
rect 11058 20304 11114 20360
rect 10966 19352 11022 19408
rect 11236 19610 11292 19612
rect 11316 19610 11372 19612
rect 11396 19610 11452 19612
rect 11476 19610 11532 19612
rect 11236 19558 11282 19610
rect 11282 19558 11292 19610
rect 11316 19558 11346 19610
rect 11346 19558 11358 19610
rect 11358 19558 11372 19610
rect 11396 19558 11410 19610
rect 11410 19558 11422 19610
rect 11422 19558 11452 19610
rect 11476 19558 11486 19610
rect 11486 19558 11532 19610
rect 11236 19556 11292 19558
rect 11316 19556 11372 19558
rect 11396 19556 11452 19558
rect 11476 19556 11532 19558
rect 11236 18522 11292 18524
rect 11316 18522 11372 18524
rect 11396 18522 11452 18524
rect 11476 18522 11532 18524
rect 11236 18470 11282 18522
rect 11282 18470 11292 18522
rect 11316 18470 11346 18522
rect 11346 18470 11358 18522
rect 11358 18470 11372 18522
rect 11396 18470 11410 18522
rect 11410 18470 11422 18522
rect 11422 18470 11452 18522
rect 11476 18470 11486 18522
rect 11486 18470 11532 18522
rect 11236 18468 11292 18470
rect 11316 18468 11372 18470
rect 11396 18468 11452 18470
rect 11476 18468 11532 18470
rect 11426 18128 11482 18184
rect 11150 17720 11206 17776
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 11426 17040 11482 17096
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 11794 18672 11850 18728
rect 11978 20848 12034 20904
rect 11794 18536 11850 18592
rect 11794 17856 11850 17912
rect 11794 17448 11850 17504
rect 11702 17176 11758 17232
rect 11794 17040 11850 17096
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 11058 14456 11114 14512
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 10598 9968 10654 10024
rect 10322 9152 10378 9208
rect 11058 10648 11114 10704
rect 10874 9016 10930 9072
rect 11794 14184 11850 14240
rect 11702 13776 11758 13832
rect 12438 27376 12494 27432
rect 12714 27376 12770 27432
rect 12950 27770 13006 27772
rect 13030 27770 13086 27772
rect 13110 27770 13166 27772
rect 13190 27770 13246 27772
rect 12950 27718 12996 27770
rect 12996 27718 13006 27770
rect 13030 27718 13060 27770
rect 13060 27718 13072 27770
rect 13072 27718 13086 27770
rect 13110 27718 13124 27770
rect 13124 27718 13136 27770
rect 13136 27718 13166 27770
rect 13190 27718 13200 27770
rect 13200 27718 13246 27770
rect 12950 27716 13006 27718
rect 13030 27716 13086 27718
rect 13110 27716 13166 27718
rect 13190 27716 13246 27718
rect 12950 26682 13006 26684
rect 13030 26682 13086 26684
rect 13110 26682 13166 26684
rect 13190 26682 13246 26684
rect 12950 26630 12996 26682
rect 12996 26630 13006 26682
rect 13030 26630 13060 26682
rect 13060 26630 13072 26682
rect 13072 26630 13086 26682
rect 13110 26630 13124 26682
rect 13124 26630 13136 26682
rect 13136 26630 13166 26682
rect 13190 26630 13200 26682
rect 13200 26630 13246 26682
rect 12950 26628 13006 26630
rect 13030 26628 13086 26630
rect 13110 26628 13166 26630
rect 13190 26628 13246 26630
rect 13542 30504 13598 30560
rect 13818 31884 13874 31920
rect 13818 31864 13820 31884
rect 13820 31864 13872 31884
rect 13872 31864 13874 31884
rect 14186 32680 14242 32736
rect 14002 32272 14058 32328
rect 13818 29144 13874 29200
rect 13634 27920 13690 27976
rect 12162 22072 12218 22128
rect 12254 21120 12310 21176
rect 12950 25594 13006 25596
rect 13030 25594 13086 25596
rect 13110 25594 13166 25596
rect 13190 25594 13246 25596
rect 12950 25542 12996 25594
rect 12996 25542 13006 25594
rect 13030 25542 13060 25594
rect 13060 25542 13072 25594
rect 13072 25542 13086 25594
rect 13110 25542 13124 25594
rect 13124 25542 13136 25594
rect 13136 25542 13166 25594
rect 13190 25542 13200 25594
rect 13200 25542 13246 25594
rect 12950 25540 13006 25542
rect 13030 25540 13086 25542
rect 13110 25540 13166 25542
rect 13190 25540 13246 25542
rect 13174 24656 13230 24712
rect 12950 24506 13006 24508
rect 13030 24506 13086 24508
rect 13110 24506 13166 24508
rect 13190 24506 13246 24508
rect 12950 24454 12996 24506
rect 12996 24454 13006 24506
rect 13030 24454 13060 24506
rect 13060 24454 13072 24506
rect 13072 24454 13086 24506
rect 13110 24454 13124 24506
rect 13124 24454 13136 24506
rect 13136 24454 13166 24506
rect 13190 24454 13200 24506
rect 13200 24454 13246 24506
rect 12950 24452 13006 24454
rect 13030 24452 13086 24454
rect 13110 24452 13166 24454
rect 13190 24452 13246 24454
rect 12622 23060 12624 23080
rect 12624 23060 12676 23080
rect 12676 23060 12678 23080
rect 12622 23024 12678 23060
rect 12950 23418 13006 23420
rect 13030 23418 13086 23420
rect 13110 23418 13166 23420
rect 13190 23418 13246 23420
rect 12950 23366 12996 23418
rect 12996 23366 13006 23418
rect 13030 23366 13060 23418
rect 13060 23366 13072 23418
rect 13072 23366 13086 23418
rect 13110 23366 13124 23418
rect 13124 23366 13136 23418
rect 13136 23366 13166 23418
rect 13190 23366 13200 23418
rect 13200 23366 13246 23418
rect 12950 23364 13006 23366
rect 13030 23364 13086 23366
rect 13110 23364 13166 23366
rect 13190 23364 13246 23366
rect 12950 22330 13006 22332
rect 13030 22330 13086 22332
rect 13110 22330 13166 22332
rect 13190 22330 13246 22332
rect 12950 22278 12996 22330
rect 12996 22278 13006 22330
rect 13030 22278 13060 22330
rect 13060 22278 13072 22330
rect 13072 22278 13086 22330
rect 13110 22278 13124 22330
rect 13124 22278 13136 22330
rect 13136 22278 13166 22330
rect 13190 22278 13200 22330
rect 13200 22278 13246 22330
rect 12950 22276 13006 22278
rect 13030 22276 13086 22278
rect 13110 22276 13166 22278
rect 13190 22276 13246 22278
rect 12162 20984 12218 21040
rect 12070 16904 12126 16960
rect 11978 15020 12034 15056
rect 11978 15000 11980 15020
rect 11980 15000 12032 15020
rect 12032 15000 12034 15020
rect 11978 14728 12034 14784
rect 11978 14476 12034 14512
rect 11978 14456 11980 14476
rect 11980 14456 12032 14476
rect 12032 14456 12034 14476
rect 12346 20304 12402 20360
rect 12806 21528 12862 21584
rect 12950 21242 13006 21244
rect 13030 21242 13086 21244
rect 13110 21242 13166 21244
rect 13190 21242 13246 21244
rect 12950 21190 12996 21242
rect 12996 21190 13006 21242
rect 13030 21190 13060 21242
rect 13060 21190 13072 21242
rect 13072 21190 13086 21242
rect 13110 21190 13124 21242
rect 13124 21190 13136 21242
rect 13136 21190 13166 21242
rect 13190 21190 13200 21242
rect 13200 21190 13246 21242
rect 12950 21188 13006 21190
rect 13030 21188 13086 21190
rect 13110 21188 13166 21190
rect 13190 21188 13246 21190
rect 12530 20440 12586 20496
rect 12950 20154 13006 20156
rect 13030 20154 13086 20156
rect 13110 20154 13166 20156
rect 13190 20154 13246 20156
rect 12950 20102 12996 20154
rect 12996 20102 13006 20154
rect 13030 20102 13060 20154
rect 13060 20102 13072 20154
rect 13072 20102 13086 20154
rect 13110 20102 13124 20154
rect 13124 20102 13136 20154
rect 13136 20102 13166 20154
rect 13190 20102 13200 20154
rect 13200 20102 13246 20154
rect 12950 20100 13006 20102
rect 13030 20100 13086 20102
rect 13110 20100 13166 20102
rect 13190 20100 13246 20102
rect 13082 19896 13138 19952
rect 13818 28464 13874 28520
rect 13818 27376 13874 27432
rect 14663 34842 14719 34844
rect 14743 34842 14799 34844
rect 14823 34842 14879 34844
rect 14903 34842 14959 34844
rect 14663 34790 14709 34842
rect 14709 34790 14719 34842
rect 14743 34790 14773 34842
rect 14773 34790 14785 34842
rect 14785 34790 14799 34842
rect 14823 34790 14837 34842
rect 14837 34790 14849 34842
rect 14849 34790 14879 34842
rect 14903 34790 14913 34842
rect 14913 34790 14959 34842
rect 14663 34788 14719 34790
rect 14743 34788 14799 34790
rect 14823 34788 14879 34790
rect 14903 34788 14959 34790
rect 14554 33904 14610 33960
rect 14663 33754 14719 33756
rect 14743 33754 14799 33756
rect 14823 33754 14879 33756
rect 14903 33754 14959 33756
rect 14663 33702 14709 33754
rect 14709 33702 14719 33754
rect 14743 33702 14773 33754
rect 14773 33702 14785 33754
rect 14785 33702 14799 33754
rect 14823 33702 14837 33754
rect 14837 33702 14849 33754
rect 14849 33702 14879 33754
rect 14903 33702 14913 33754
rect 14913 33702 14959 33754
rect 14663 33700 14719 33702
rect 14743 33700 14799 33702
rect 14823 33700 14879 33702
rect 14903 33700 14959 33702
rect 14278 30640 14334 30696
rect 14278 28600 14334 28656
rect 14186 26968 14242 27024
rect 13634 25780 13636 25800
rect 13636 25780 13688 25800
rect 13688 25780 13690 25800
rect 13634 25744 13690 25780
rect 13542 22480 13598 22536
rect 14002 24656 14058 24712
rect 13910 24112 13966 24168
rect 14186 25644 14188 25664
rect 14188 25644 14240 25664
rect 14240 25644 14242 25664
rect 14186 25608 14242 25644
rect 12438 17992 12494 18048
rect 12530 17312 12586 17368
rect 12950 19066 13006 19068
rect 13030 19066 13086 19068
rect 13110 19066 13166 19068
rect 13190 19066 13246 19068
rect 12950 19014 12996 19066
rect 12996 19014 13006 19066
rect 13030 19014 13060 19066
rect 13060 19014 13072 19066
rect 13072 19014 13086 19066
rect 13110 19014 13124 19066
rect 13124 19014 13136 19066
rect 13136 19014 13166 19066
rect 13190 19014 13200 19066
rect 13200 19014 13246 19066
rect 12950 19012 13006 19014
rect 13030 19012 13086 19014
rect 13110 19012 13166 19014
rect 13190 19012 13246 19014
rect 12990 18808 13046 18864
rect 12530 16788 12586 16824
rect 12530 16768 12532 16788
rect 12532 16768 12584 16788
rect 12584 16768 12586 16788
rect 12950 17978 13006 17980
rect 13030 17978 13086 17980
rect 13110 17978 13166 17980
rect 13190 17978 13246 17980
rect 12950 17926 12996 17978
rect 12996 17926 13006 17978
rect 13030 17926 13060 17978
rect 13060 17926 13072 17978
rect 13072 17926 13086 17978
rect 13110 17926 13124 17978
rect 13124 17926 13136 17978
rect 13136 17926 13166 17978
rect 13190 17926 13200 17978
rect 13200 17926 13246 17978
rect 12950 17924 13006 17926
rect 13030 17924 13086 17926
rect 13110 17924 13166 17926
rect 13190 17924 13246 17926
rect 13726 22344 13782 22400
rect 13818 22072 13874 22128
rect 13634 21528 13690 21584
rect 14186 23468 14188 23488
rect 14188 23468 14240 23488
rect 14240 23468 14242 23488
rect 14186 23432 14242 23468
rect 13910 20984 13966 21040
rect 13910 19896 13966 19952
rect 13818 19352 13874 19408
rect 14094 21528 14150 21584
rect 14094 18808 14150 18864
rect 13910 18536 13966 18592
rect 13910 18264 13966 18320
rect 13818 17876 13874 17912
rect 13818 17856 13820 17876
rect 13820 17856 13872 17876
rect 13872 17856 13874 17876
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 12898 16632 12954 16688
rect 12714 14728 12770 14784
rect 12254 13232 12310 13288
rect 11794 12280 11850 12336
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 11702 10920 11758 10976
rect 11886 11212 11942 11248
rect 11886 11192 11888 11212
rect 11888 11192 11940 11212
rect 11940 11192 11942 11212
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 11242 9288 11298 9344
rect 11426 9016 11482 9072
rect 11150 8880 11206 8936
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 11886 9424 11942 9480
rect 11794 9288 11850 9344
rect 11702 9152 11758 9208
rect 11518 8472 11574 8528
rect 11978 9016 12034 9072
rect 11978 8880 12034 8936
rect 11334 7792 11390 7848
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 12254 12844 12310 12880
rect 12254 12824 12256 12844
rect 12256 12824 12308 12844
rect 12308 12824 12310 12844
rect 12530 13912 12586 13968
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 13266 15544 13322 15600
rect 13082 15136 13138 15192
rect 12990 14864 13046 14920
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 12622 13232 12678 13288
rect 12254 9696 12310 9752
rect 12162 9560 12218 9616
rect 12714 10124 12770 10160
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 13266 12180 13268 12200
rect 13268 12180 13320 12200
rect 13320 12180 13322 12200
rect 13266 12144 13322 12180
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 12714 10104 12716 10124
rect 12716 10104 12768 10124
rect 12768 10104 12770 10124
rect 12806 9968 12862 10024
rect 12346 9152 12402 9208
rect 12714 8608 12770 8664
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 12162 7792 12218 7848
rect 12346 6840 12402 6896
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 12438 6316 12494 6352
rect 12438 6296 12440 6316
rect 12440 6296 12492 6316
rect 12492 6296 12494 6316
rect 12806 8336 12862 8392
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 13726 17448 13782 17504
rect 13450 15952 13506 16008
rect 13726 16360 13782 16416
rect 14370 23160 14426 23216
rect 14278 22616 14334 22672
rect 14663 32666 14719 32668
rect 14743 32666 14799 32668
rect 14823 32666 14879 32668
rect 14903 32666 14959 32668
rect 14663 32614 14709 32666
rect 14709 32614 14719 32666
rect 14743 32614 14773 32666
rect 14773 32614 14785 32666
rect 14785 32614 14799 32666
rect 14823 32614 14837 32666
rect 14837 32614 14849 32666
rect 14849 32614 14879 32666
rect 14903 32614 14913 32666
rect 14913 32614 14959 32666
rect 14663 32612 14719 32614
rect 14743 32612 14799 32614
rect 14823 32612 14879 32614
rect 14903 32612 14959 32614
rect 14663 31578 14719 31580
rect 14743 31578 14799 31580
rect 14823 31578 14879 31580
rect 14903 31578 14959 31580
rect 14663 31526 14709 31578
rect 14709 31526 14719 31578
rect 14743 31526 14773 31578
rect 14773 31526 14785 31578
rect 14785 31526 14799 31578
rect 14823 31526 14837 31578
rect 14837 31526 14849 31578
rect 14849 31526 14879 31578
rect 14903 31526 14913 31578
rect 14913 31526 14959 31578
rect 14663 31524 14719 31526
rect 14743 31524 14799 31526
rect 14823 31524 14879 31526
rect 14903 31524 14959 31526
rect 14554 30776 14610 30832
rect 14663 30490 14719 30492
rect 14743 30490 14799 30492
rect 14823 30490 14879 30492
rect 14903 30490 14959 30492
rect 14663 30438 14709 30490
rect 14709 30438 14719 30490
rect 14743 30438 14773 30490
rect 14773 30438 14785 30490
rect 14785 30438 14799 30490
rect 14823 30438 14837 30490
rect 14837 30438 14849 30490
rect 14849 30438 14879 30490
rect 14903 30438 14913 30490
rect 14913 30438 14959 30490
rect 14663 30436 14719 30438
rect 14743 30436 14799 30438
rect 14823 30436 14879 30438
rect 14903 30436 14959 30438
rect 14663 29402 14719 29404
rect 14743 29402 14799 29404
rect 14823 29402 14879 29404
rect 14903 29402 14959 29404
rect 14663 29350 14709 29402
rect 14709 29350 14719 29402
rect 14743 29350 14773 29402
rect 14773 29350 14785 29402
rect 14785 29350 14799 29402
rect 14823 29350 14837 29402
rect 14837 29350 14849 29402
rect 14849 29350 14879 29402
rect 14903 29350 14913 29402
rect 14913 29350 14959 29402
rect 14663 29348 14719 29350
rect 14743 29348 14799 29350
rect 14823 29348 14879 29350
rect 14903 29348 14959 29350
rect 14663 28314 14719 28316
rect 14743 28314 14799 28316
rect 14823 28314 14879 28316
rect 14903 28314 14959 28316
rect 14663 28262 14709 28314
rect 14709 28262 14719 28314
rect 14743 28262 14773 28314
rect 14773 28262 14785 28314
rect 14785 28262 14799 28314
rect 14823 28262 14837 28314
rect 14837 28262 14849 28314
rect 14849 28262 14879 28314
rect 14903 28262 14913 28314
rect 14913 28262 14959 28314
rect 14663 28260 14719 28262
rect 14743 28260 14799 28262
rect 14823 28260 14879 28262
rect 14903 28260 14959 28262
rect 14663 27226 14719 27228
rect 14743 27226 14799 27228
rect 14823 27226 14879 27228
rect 14903 27226 14959 27228
rect 14663 27174 14709 27226
rect 14709 27174 14719 27226
rect 14743 27174 14773 27226
rect 14773 27174 14785 27226
rect 14785 27174 14799 27226
rect 14823 27174 14837 27226
rect 14837 27174 14849 27226
rect 14849 27174 14879 27226
rect 14903 27174 14913 27226
rect 14913 27174 14959 27226
rect 14663 27172 14719 27174
rect 14743 27172 14799 27174
rect 14823 27172 14879 27174
rect 14903 27172 14959 27174
rect 14646 26696 14702 26752
rect 14663 26138 14719 26140
rect 14743 26138 14799 26140
rect 14823 26138 14879 26140
rect 14903 26138 14959 26140
rect 14663 26086 14709 26138
rect 14709 26086 14719 26138
rect 14743 26086 14773 26138
rect 14773 26086 14785 26138
rect 14785 26086 14799 26138
rect 14823 26086 14837 26138
rect 14837 26086 14849 26138
rect 14849 26086 14879 26138
rect 14903 26086 14913 26138
rect 14913 26086 14959 26138
rect 14663 26084 14719 26086
rect 14743 26084 14799 26086
rect 14823 26084 14879 26086
rect 14903 26084 14959 26086
rect 14554 25472 14610 25528
rect 14370 21936 14426 21992
rect 14278 20984 14334 21040
rect 14370 20168 14426 20224
rect 14278 19080 14334 19136
rect 14186 17448 14242 17504
rect 14663 25050 14719 25052
rect 14743 25050 14799 25052
rect 14823 25050 14879 25052
rect 14903 25050 14959 25052
rect 14663 24998 14709 25050
rect 14709 24998 14719 25050
rect 14743 24998 14773 25050
rect 14773 24998 14785 25050
rect 14785 24998 14799 25050
rect 14823 24998 14837 25050
rect 14837 24998 14849 25050
rect 14849 24998 14879 25050
rect 14903 24998 14913 25050
rect 14913 24998 14959 25050
rect 14663 24996 14719 24998
rect 14743 24996 14799 24998
rect 14823 24996 14879 24998
rect 14903 24996 14959 24998
rect 14663 23962 14719 23964
rect 14743 23962 14799 23964
rect 14823 23962 14879 23964
rect 14903 23962 14959 23964
rect 14663 23910 14709 23962
rect 14709 23910 14719 23962
rect 14743 23910 14773 23962
rect 14773 23910 14785 23962
rect 14785 23910 14799 23962
rect 14823 23910 14837 23962
rect 14837 23910 14849 23962
rect 14849 23910 14879 23962
rect 14903 23910 14913 23962
rect 14913 23910 14959 23962
rect 14663 23908 14719 23910
rect 14743 23908 14799 23910
rect 14823 23908 14879 23910
rect 14903 23908 14959 23910
rect 14663 22874 14719 22876
rect 14743 22874 14799 22876
rect 14823 22874 14879 22876
rect 14903 22874 14959 22876
rect 14663 22822 14709 22874
rect 14709 22822 14719 22874
rect 14743 22822 14773 22874
rect 14773 22822 14785 22874
rect 14785 22822 14799 22874
rect 14823 22822 14837 22874
rect 14837 22822 14849 22874
rect 14849 22822 14879 22874
rect 14903 22822 14913 22874
rect 14913 22822 14959 22874
rect 14663 22820 14719 22822
rect 14743 22820 14799 22822
rect 14823 22820 14879 22822
rect 14903 22820 14959 22822
rect 14663 21786 14719 21788
rect 14743 21786 14799 21788
rect 14823 21786 14879 21788
rect 14903 21786 14959 21788
rect 14663 21734 14709 21786
rect 14709 21734 14719 21786
rect 14743 21734 14773 21786
rect 14773 21734 14785 21786
rect 14785 21734 14799 21786
rect 14823 21734 14837 21786
rect 14837 21734 14849 21786
rect 14849 21734 14879 21786
rect 14903 21734 14913 21786
rect 14913 21734 14959 21786
rect 14663 21732 14719 21734
rect 14743 21732 14799 21734
rect 14823 21732 14879 21734
rect 14903 21732 14959 21734
rect 14663 20698 14719 20700
rect 14743 20698 14799 20700
rect 14823 20698 14879 20700
rect 14903 20698 14959 20700
rect 14663 20646 14709 20698
rect 14709 20646 14719 20698
rect 14743 20646 14773 20698
rect 14773 20646 14785 20698
rect 14785 20646 14799 20698
rect 14823 20646 14837 20698
rect 14837 20646 14849 20698
rect 14849 20646 14879 20698
rect 14903 20646 14913 20698
rect 14913 20646 14959 20698
rect 14663 20644 14719 20646
rect 14743 20644 14799 20646
rect 14823 20644 14879 20646
rect 14903 20644 14959 20646
rect 14663 19610 14719 19612
rect 14743 19610 14799 19612
rect 14823 19610 14879 19612
rect 14903 19610 14959 19612
rect 14663 19558 14709 19610
rect 14709 19558 14719 19610
rect 14743 19558 14773 19610
rect 14773 19558 14785 19610
rect 14785 19558 14799 19610
rect 14823 19558 14837 19610
rect 14837 19558 14849 19610
rect 14849 19558 14879 19610
rect 14903 19558 14913 19610
rect 14913 19558 14959 19610
rect 14663 19556 14719 19558
rect 14743 19556 14799 19558
rect 14823 19556 14879 19558
rect 14903 19556 14959 19558
rect 14663 18522 14719 18524
rect 14743 18522 14799 18524
rect 14823 18522 14879 18524
rect 14903 18522 14959 18524
rect 14663 18470 14709 18522
rect 14709 18470 14719 18522
rect 14743 18470 14773 18522
rect 14773 18470 14785 18522
rect 14785 18470 14799 18522
rect 14823 18470 14837 18522
rect 14837 18470 14849 18522
rect 14849 18470 14879 18522
rect 14903 18470 14913 18522
rect 14913 18470 14959 18522
rect 14663 18468 14719 18470
rect 14743 18468 14799 18470
rect 14823 18468 14879 18470
rect 14903 18468 14959 18470
rect 14278 16632 14334 16688
rect 14186 16360 14242 16416
rect 14186 16088 14242 16144
rect 13726 13912 13782 13968
rect 14094 15408 14150 15464
rect 14094 15272 14150 15328
rect 14278 14728 14334 14784
rect 14186 13776 14242 13832
rect 13910 12824 13966 12880
rect 13910 12552 13966 12608
rect 13726 11872 13782 11928
rect 13634 10512 13690 10568
rect 13450 9424 13506 9480
rect 13910 11736 13966 11792
rect 13910 10104 13966 10160
rect 13818 9288 13874 9344
rect 13358 7928 13414 7984
rect 13726 7384 13782 7440
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 12898 6296 12954 6352
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 13358 5752 13414 5808
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 12438 3440 12494 3496
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 11058 2624 11114 2680
rect 9523 1658 9579 1660
rect 9603 1658 9659 1660
rect 9683 1658 9739 1660
rect 9763 1658 9819 1660
rect 9523 1606 9569 1658
rect 9569 1606 9579 1658
rect 9603 1606 9633 1658
rect 9633 1606 9645 1658
rect 9645 1606 9659 1658
rect 9683 1606 9697 1658
rect 9697 1606 9709 1658
rect 9709 1606 9739 1658
rect 9763 1606 9773 1658
rect 9773 1606 9819 1658
rect 9523 1604 9579 1606
rect 9603 1604 9659 1606
rect 9683 1604 9739 1606
rect 9763 1604 9819 1606
rect 11794 2624 11850 2680
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 13726 7112 13782 7168
rect 13634 6724 13690 6760
rect 13634 6704 13636 6724
rect 13636 6704 13688 6724
rect 13688 6704 13690 6724
rect 13726 5208 13782 5264
rect 13910 6196 13912 6216
rect 13912 6196 13964 6216
rect 13964 6196 13966 6216
rect 13910 6160 13966 6196
rect 13910 5616 13966 5672
rect 14186 13368 14242 13424
rect 14554 17856 14610 17912
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 14554 17040 14610 17096
rect 14554 16904 14610 16960
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 14278 12824 14334 12880
rect 14278 12008 14334 12064
rect 14186 11736 14242 11792
rect 14186 10376 14242 10432
rect 14278 9560 14334 9616
rect 14278 8200 14334 8256
rect 14186 6024 14242 6080
rect 14462 12708 14518 12744
rect 14462 12688 14464 12708
rect 14464 12688 14516 12708
rect 14516 12688 14518 12708
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 14646 13640 14702 13696
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 14646 11464 14702 11520
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 14186 5616 14242 5672
rect 14738 6316 14794 6352
rect 14738 6296 14740 6316
rect 14740 6296 14792 6316
rect 14792 6296 14794 6316
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 15106 37168 15162 37224
rect 15106 35980 15108 36000
rect 15108 35980 15160 36000
rect 15160 35980 15162 36000
rect 15106 35944 15162 35980
rect 15106 34856 15162 34912
rect 15106 26152 15162 26208
rect 15106 23976 15162 24032
rect 15106 22924 15108 22944
rect 15108 22924 15160 22944
rect 15160 22924 15162 22944
rect 15106 22888 15162 22924
rect 15382 35808 15438 35864
rect 15382 34448 15438 34504
rect 15382 33904 15438 33960
rect 15566 34448 15622 34504
rect 15566 32136 15622 32192
rect 15474 31592 15530 31648
rect 15658 30504 15714 30560
rect 15566 28328 15622 28384
rect 15474 27512 15530 27568
rect 15474 25880 15530 25936
rect 15198 21800 15254 21856
rect 15198 17856 15254 17912
rect 15198 17448 15254 17504
rect 15198 13096 15254 13152
rect 15106 12008 15162 12064
rect 15106 10104 15162 10160
rect 15106 7656 15162 7712
rect 15106 6568 15162 6624
rect 15106 5480 15162 5536
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
rect 12950 1658 13006 1660
rect 13030 1658 13086 1660
rect 13110 1658 13166 1660
rect 13190 1658 13246 1660
rect 12950 1606 12996 1658
rect 12996 1606 13006 1658
rect 13030 1606 13060 1658
rect 13060 1606 13072 1658
rect 13072 1606 13086 1658
rect 13110 1606 13124 1658
rect 13124 1606 13136 1658
rect 13136 1606 13166 1658
rect 13190 1606 13200 1658
rect 13200 1606 13246 1658
rect 12950 1604 13006 1606
rect 13030 1604 13086 1606
rect 13110 1604 13166 1606
rect 13190 1604 13246 1606
rect 15474 19624 15530 19680
rect 15474 14456 15530 14512
rect 15474 14048 15530 14104
rect 15658 15816 15714 15872
rect 15474 9832 15530 9888
rect 4618 1300 4620 1320
rect 4620 1300 4672 1320
rect 4672 1300 4674 1320
rect 4618 1264 4674 1300
rect 5354 1300 5356 1320
rect 5356 1300 5408 1320
rect 5408 1300 5410 1320
rect 5354 1264 5410 1300
rect 4382 1114 4438 1116
rect 4462 1114 4518 1116
rect 4542 1114 4598 1116
rect 4622 1114 4678 1116
rect 4382 1062 4428 1114
rect 4428 1062 4438 1114
rect 4462 1062 4492 1114
rect 4492 1062 4504 1114
rect 4504 1062 4518 1114
rect 4542 1062 4556 1114
rect 4556 1062 4568 1114
rect 4568 1062 4598 1114
rect 4622 1062 4632 1114
rect 4632 1062 4678 1114
rect 4382 1060 4438 1062
rect 4462 1060 4518 1062
rect 4542 1060 4598 1062
rect 4622 1060 4678 1062
rect 7809 1114 7865 1116
rect 7889 1114 7945 1116
rect 7969 1114 8025 1116
rect 8049 1114 8105 1116
rect 7809 1062 7855 1114
rect 7855 1062 7865 1114
rect 7889 1062 7919 1114
rect 7919 1062 7931 1114
rect 7931 1062 7945 1114
rect 7969 1062 7983 1114
rect 7983 1062 7995 1114
rect 7995 1062 8025 1114
rect 8049 1062 8059 1114
rect 8059 1062 8105 1114
rect 7809 1060 7865 1062
rect 7889 1060 7945 1062
rect 7969 1060 8025 1062
rect 8049 1060 8105 1062
rect 11236 1114 11292 1116
rect 11316 1114 11372 1116
rect 11396 1114 11452 1116
rect 11476 1114 11532 1116
rect 11236 1062 11282 1114
rect 11282 1062 11292 1114
rect 11316 1062 11346 1114
rect 11346 1062 11358 1114
rect 11358 1062 11372 1114
rect 11396 1062 11410 1114
rect 11410 1062 11422 1114
rect 11422 1062 11452 1114
rect 11476 1062 11486 1114
rect 11486 1062 11532 1114
rect 11236 1060 11292 1062
rect 11316 1060 11372 1062
rect 11396 1060 11452 1062
rect 11476 1060 11532 1062
rect 14663 1114 14719 1116
rect 14743 1114 14799 1116
rect 14823 1114 14879 1116
rect 14903 1114 14959 1116
rect 14663 1062 14709 1114
rect 14709 1062 14719 1114
rect 14743 1062 14773 1114
rect 14773 1062 14785 1114
rect 14785 1062 14799 1114
rect 14823 1062 14837 1114
rect 14837 1062 14849 1114
rect 14849 1062 14879 1114
rect 14903 1062 14913 1114
rect 14913 1062 14959 1114
rect 14663 1060 14719 1062
rect 14743 1060 14799 1062
rect 14823 1060 14879 1062
rect 14903 1060 14959 1062
<< metal3 >>
rect 4372 43552 4688 43553
rect 4372 43488 4378 43552
rect 4442 43488 4458 43552
rect 4522 43488 4538 43552
rect 4602 43488 4618 43552
rect 4682 43488 4688 43552
rect 4372 43487 4688 43488
rect 7799 43552 8115 43553
rect 7799 43488 7805 43552
rect 7869 43488 7885 43552
rect 7949 43488 7965 43552
rect 8029 43488 8045 43552
rect 8109 43488 8115 43552
rect 7799 43487 8115 43488
rect 11226 43552 11542 43553
rect 11226 43488 11232 43552
rect 11296 43488 11312 43552
rect 11376 43488 11392 43552
rect 11456 43488 11472 43552
rect 11536 43488 11542 43552
rect 11226 43487 11542 43488
rect 14653 43552 14969 43553
rect 14653 43488 14659 43552
rect 14723 43488 14739 43552
rect 14803 43488 14819 43552
rect 14883 43488 14899 43552
rect 14963 43488 14969 43552
rect 14653 43487 14969 43488
rect 2659 43008 2975 43009
rect 2659 42944 2665 43008
rect 2729 42944 2745 43008
rect 2809 42944 2825 43008
rect 2889 42944 2905 43008
rect 2969 42944 2975 43008
rect 2659 42943 2975 42944
rect 6086 43008 6402 43009
rect 6086 42944 6092 43008
rect 6156 42944 6172 43008
rect 6236 42944 6252 43008
rect 6316 42944 6332 43008
rect 6396 42944 6402 43008
rect 6086 42943 6402 42944
rect 9513 43008 9829 43009
rect 9513 42944 9519 43008
rect 9583 42944 9599 43008
rect 9663 42944 9679 43008
rect 9743 42944 9759 43008
rect 9823 42944 9829 43008
rect 9513 42943 9829 42944
rect 12940 43008 13256 43009
rect 12940 42944 12946 43008
rect 13010 42944 13026 43008
rect 13090 42944 13106 43008
rect 13170 42944 13186 43008
rect 13250 42944 13256 43008
rect 12940 42943 13256 42944
rect 6678 42604 6684 42668
rect 6748 42666 6754 42668
rect 12433 42666 12499 42669
rect 6748 42664 12499 42666
rect 6748 42608 12438 42664
rect 12494 42608 12499 42664
rect 6748 42606 12499 42608
rect 6748 42604 6754 42606
rect 12433 42603 12499 42606
rect 4372 42464 4688 42465
rect 4372 42400 4378 42464
rect 4442 42400 4458 42464
rect 4522 42400 4538 42464
rect 4602 42400 4618 42464
rect 4682 42400 4688 42464
rect 4372 42399 4688 42400
rect 7799 42464 8115 42465
rect 7799 42400 7805 42464
rect 7869 42400 7885 42464
rect 7949 42400 7965 42464
rect 8029 42400 8045 42464
rect 8109 42400 8115 42464
rect 7799 42399 8115 42400
rect 11226 42464 11542 42465
rect 11226 42400 11232 42464
rect 11296 42400 11312 42464
rect 11376 42400 11392 42464
rect 11456 42400 11472 42464
rect 11536 42400 11542 42464
rect 11226 42399 11542 42400
rect 14653 42464 14969 42465
rect 14653 42400 14659 42464
rect 14723 42400 14739 42464
rect 14803 42400 14819 42464
rect 14883 42400 14899 42464
rect 14963 42400 14969 42464
rect 14653 42399 14969 42400
rect 2659 41920 2975 41921
rect 2659 41856 2665 41920
rect 2729 41856 2745 41920
rect 2809 41856 2825 41920
rect 2889 41856 2905 41920
rect 2969 41856 2975 41920
rect 2659 41855 2975 41856
rect 6086 41920 6402 41921
rect 6086 41856 6092 41920
rect 6156 41856 6172 41920
rect 6236 41856 6252 41920
rect 6316 41856 6332 41920
rect 6396 41856 6402 41920
rect 6086 41855 6402 41856
rect 9513 41920 9829 41921
rect 9513 41856 9519 41920
rect 9583 41856 9599 41920
rect 9663 41856 9679 41920
rect 9743 41856 9759 41920
rect 9823 41856 9829 41920
rect 9513 41855 9829 41856
rect 12940 41920 13256 41921
rect 12940 41856 12946 41920
rect 13010 41856 13026 41920
rect 13090 41856 13106 41920
rect 13170 41856 13186 41920
rect 13250 41856 13256 41920
rect 12940 41855 13256 41856
rect 2262 41652 2268 41716
rect 2332 41714 2338 41716
rect 9397 41714 9463 41717
rect 2332 41712 9463 41714
rect 2332 41656 9402 41712
rect 9458 41656 9463 41712
rect 2332 41654 9463 41656
rect 2332 41652 2338 41654
rect 9397 41651 9463 41654
rect 4245 41578 4311 41581
rect 4838 41578 4844 41580
rect 4245 41576 4844 41578
rect 4245 41520 4250 41576
rect 4306 41520 4844 41576
rect 4245 41518 4844 41520
rect 4245 41515 4311 41518
rect 4838 41516 4844 41518
rect 4908 41516 4914 41580
rect 7414 41516 7420 41580
rect 7484 41578 7490 41580
rect 11697 41578 11763 41581
rect 7484 41576 11763 41578
rect 7484 41520 11702 41576
rect 11758 41520 11763 41576
rect 7484 41518 11763 41520
rect 7484 41516 7490 41518
rect 11697 41515 11763 41518
rect 5073 41442 5139 41445
rect 10961 41444 11027 41445
rect 5390 41442 5396 41444
rect 5073 41440 5396 41442
rect 5073 41384 5078 41440
rect 5134 41384 5396 41440
rect 5073 41382 5396 41384
rect 5073 41379 5139 41382
rect 5390 41380 5396 41382
rect 5460 41380 5466 41444
rect 10910 41442 10916 41444
rect 10870 41382 10916 41442
rect 10980 41440 11027 41444
rect 11022 41384 11027 41440
rect 10910 41380 10916 41382
rect 10980 41380 11027 41384
rect 10961 41379 11027 41380
rect 4372 41376 4688 41377
rect 4372 41312 4378 41376
rect 4442 41312 4458 41376
rect 4522 41312 4538 41376
rect 4602 41312 4618 41376
rect 4682 41312 4688 41376
rect 4372 41311 4688 41312
rect 7799 41376 8115 41377
rect 7799 41312 7805 41376
rect 7869 41312 7885 41376
rect 7949 41312 7965 41376
rect 8029 41312 8045 41376
rect 8109 41312 8115 41376
rect 7799 41311 8115 41312
rect 11226 41376 11542 41377
rect 11226 41312 11232 41376
rect 11296 41312 11312 41376
rect 11376 41312 11392 41376
rect 11456 41312 11472 41376
rect 11536 41312 11542 41376
rect 11226 41311 11542 41312
rect 14653 41376 14969 41377
rect 14653 41312 14659 41376
rect 14723 41312 14739 41376
rect 14803 41312 14819 41376
rect 14883 41312 14899 41376
rect 14963 41312 14969 41376
rect 14653 41311 14969 41312
rect 0 40898 160 40928
rect 749 40898 815 40901
rect 0 40896 815 40898
rect 0 40840 754 40896
rect 810 40840 815 40896
rect 0 40838 815 40840
rect 0 40808 160 40838
rect 749 40835 815 40838
rect 2659 40832 2975 40833
rect 2659 40768 2665 40832
rect 2729 40768 2745 40832
rect 2809 40768 2825 40832
rect 2889 40768 2905 40832
rect 2969 40768 2975 40832
rect 2659 40767 2975 40768
rect 6086 40832 6402 40833
rect 6086 40768 6092 40832
rect 6156 40768 6172 40832
rect 6236 40768 6252 40832
rect 6316 40768 6332 40832
rect 6396 40768 6402 40832
rect 6086 40767 6402 40768
rect 9513 40832 9829 40833
rect 9513 40768 9519 40832
rect 9583 40768 9599 40832
rect 9663 40768 9679 40832
rect 9743 40768 9759 40832
rect 9823 40768 9829 40832
rect 9513 40767 9829 40768
rect 12940 40832 13256 40833
rect 12940 40768 12946 40832
rect 13010 40768 13026 40832
rect 13090 40768 13106 40832
rect 13170 40768 13186 40832
rect 13250 40768 13256 40832
rect 12940 40767 13256 40768
rect 4372 40288 4688 40289
rect 4372 40224 4378 40288
rect 4442 40224 4458 40288
rect 4522 40224 4538 40288
rect 4602 40224 4618 40288
rect 4682 40224 4688 40288
rect 4372 40223 4688 40224
rect 7799 40288 8115 40289
rect 7799 40224 7805 40288
rect 7869 40224 7885 40288
rect 7949 40224 7965 40288
rect 8029 40224 8045 40288
rect 8109 40224 8115 40288
rect 7799 40223 8115 40224
rect 11226 40288 11542 40289
rect 11226 40224 11232 40288
rect 11296 40224 11312 40288
rect 11376 40224 11392 40288
rect 11456 40224 11472 40288
rect 11536 40224 11542 40288
rect 11226 40223 11542 40224
rect 14653 40288 14969 40289
rect 14653 40224 14659 40288
rect 14723 40224 14739 40288
rect 14803 40224 14819 40288
rect 14883 40224 14899 40288
rect 14963 40224 14969 40288
rect 14653 40223 14969 40224
rect 0 40082 160 40112
rect 749 40082 815 40085
rect 9305 40084 9371 40085
rect 0 40080 815 40082
rect 0 40024 754 40080
rect 810 40024 815 40080
rect 0 40022 815 40024
rect 0 39992 160 40022
rect 749 40019 815 40022
rect 9254 40020 9260 40084
rect 9324 40082 9371 40084
rect 9324 40080 9416 40082
rect 9366 40024 9416 40080
rect 9324 40022 9416 40024
rect 9324 40020 9371 40022
rect 9305 40019 9371 40020
rect 13721 39810 13787 39813
rect 15840 39810 16000 39840
rect 13721 39808 16000 39810
rect 13721 39752 13726 39808
rect 13782 39752 16000 39808
rect 13721 39750 16000 39752
rect 13721 39747 13787 39750
rect 2659 39744 2975 39745
rect 2659 39680 2665 39744
rect 2729 39680 2745 39744
rect 2809 39680 2825 39744
rect 2889 39680 2905 39744
rect 2969 39680 2975 39744
rect 2659 39679 2975 39680
rect 6086 39744 6402 39745
rect 6086 39680 6092 39744
rect 6156 39680 6172 39744
rect 6236 39680 6252 39744
rect 6316 39680 6332 39744
rect 6396 39680 6402 39744
rect 6086 39679 6402 39680
rect 9513 39744 9829 39745
rect 9513 39680 9519 39744
rect 9583 39680 9599 39744
rect 9663 39680 9679 39744
rect 9743 39680 9759 39744
rect 9823 39680 9829 39744
rect 9513 39679 9829 39680
rect 12940 39744 13256 39745
rect 12940 39680 12946 39744
rect 13010 39680 13026 39744
rect 13090 39680 13106 39744
rect 13170 39680 13186 39744
rect 13250 39680 13256 39744
rect 15840 39720 16000 39750
rect 12940 39679 13256 39680
rect 13997 39538 14063 39541
rect 14181 39538 14247 39541
rect 15840 39538 16000 39568
rect 13997 39536 14106 39538
rect 13997 39480 14002 39536
rect 14058 39480 14106 39536
rect 13997 39475 14106 39480
rect 14181 39536 16000 39538
rect 14181 39480 14186 39536
rect 14242 39480 16000 39536
rect 14181 39478 16000 39480
rect 14181 39475 14247 39478
rect 14046 39402 14106 39475
rect 15840 39448 16000 39478
rect 14046 39342 15210 39402
rect 0 39266 160 39296
rect 749 39266 815 39269
rect 0 39264 815 39266
rect 0 39208 754 39264
rect 810 39208 815 39264
rect 0 39206 815 39208
rect 15150 39266 15210 39342
rect 15840 39266 16000 39296
rect 15150 39206 16000 39266
rect 0 39176 160 39206
rect 749 39203 815 39206
rect 4372 39200 4688 39201
rect 4372 39136 4378 39200
rect 4442 39136 4458 39200
rect 4522 39136 4538 39200
rect 4602 39136 4618 39200
rect 4682 39136 4688 39200
rect 4372 39135 4688 39136
rect 7799 39200 8115 39201
rect 7799 39136 7805 39200
rect 7869 39136 7885 39200
rect 7949 39136 7965 39200
rect 8029 39136 8045 39200
rect 8109 39136 8115 39200
rect 7799 39135 8115 39136
rect 11226 39200 11542 39201
rect 11226 39136 11232 39200
rect 11296 39136 11312 39200
rect 11376 39136 11392 39200
rect 11456 39136 11472 39200
rect 11536 39136 11542 39200
rect 11226 39135 11542 39136
rect 14653 39200 14969 39201
rect 14653 39136 14659 39200
rect 14723 39136 14739 39200
rect 14803 39136 14819 39200
rect 14883 39136 14899 39200
rect 14963 39136 14969 39200
rect 15840 39176 16000 39206
rect 14653 39135 14969 39136
rect 13905 38994 13971 38997
rect 15840 38994 16000 39024
rect 13905 38992 16000 38994
rect 13905 38936 13910 38992
rect 13966 38936 16000 38992
rect 13905 38934 16000 38936
rect 13905 38931 13971 38934
rect 15840 38904 16000 38934
rect 14365 38722 14431 38725
rect 15840 38722 16000 38752
rect 14365 38720 16000 38722
rect 14365 38664 14370 38720
rect 14426 38664 16000 38720
rect 14365 38662 16000 38664
rect 14365 38659 14431 38662
rect 2659 38656 2975 38657
rect 2659 38592 2665 38656
rect 2729 38592 2745 38656
rect 2809 38592 2825 38656
rect 2889 38592 2905 38656
rect 2969 38592 2975 38656
rect 2659 38591 2975 38592
rect 6086 38656 6402 38657
rect 6086 38592 6092 38656
rect 6156 38592 6172 38656
rect 6236 38592 6252 38656
rect 6316 38592 6332 38656
rect 6396 38592 6402 38656
rect 6086 38591 6402 38592
rect 9513 38656 9829 38657
rect 9513 38592 9519 38656
rect 9583 38592 9599 38656
rect 9663 38592 9679 38656
rect 9743 38592 9759 38656
rect 9823 38592 9829 38656
rect 9513 38591 9829 38592
rect 12940 38656 13256 38657
rect 12940 38592 12946 38656
rect 13010 38592 13026 38656
rect 13090 38592 13106 38656
rect 13170 38592 13186 38656
rect 13250 38592 13256 38656
rect 15840 38632 16000 38662
rect 12940 38591 13256 38592
rect 1393 38586 1459 38589
rect 798 38584 1459 38586
rect 798 38528 1398 38584
rect 1454 38528 1459 38584
rect 798 38526 1459 38528
rect 0 38450 160 38480
rect 798 38450 858 38526
rect 1393 38523 1459 38526
rect 14181 38586 14247 38589
rect 14181 38584 15026 38586
rect 14181 38528 14186 38584
rect 14242 38528 15026 38584
rect 14181 38526 15026 38528
rect 14181 38523 14247 38526
rect 0 38390 858 38450
rect 13629 38450 13695 38453
rect 14966 38450 15026 38526
rect 15840 38450 16000 38480
rect 13629 38448 14842 38450
rect 13629 38392 13634 38448
rect 13690 38392 14842 38448
rect 13629 38390 14842 38392
rect 14966 38390 16000 38450
rect 0 38360 160 38390
rect 13629 38387 13695 38390
rect 14782 38314 14842 38390
rect 15840 38360 16000 38390
rect 14782 38254 15210 38314
rect 15150 38178 15210 38254
rect 15840 38178 16000 38208
rect 15150 38118 16000 38178
rect 4372 38112 4688 38113
rect 4372 38048 4378 38112
rect 4442 38048 4458 38112
rect 4522 38048 4538 38112
rect 4602 38048 4618 38112
rect 4682 38048 4688 38112
rect 4372 38047 4688 38048
rect 7799 38112 8115 38113
rect 7799 38048 7805 38112
rect 7869 38048 7885 38112
rect 7949 38048 7965 38112
rect 8029 38048 8045 38112
rect 8109 38048 8115 38112
rect 7799 38047 8115 38048
rect 11226 38112 11542 38113
rect 11226 38048 11232 38112
rect 11296 38048 11312 38112
rect 11376 38048 11392 38112
rect 11456 38048 11472 38112
rect 11536 38048 11542 38112
rect 11226 38047 11542 38048
rect 14653 38112 14969 38113
rect 14653 38048 14659 38112
rect 14723 38048 14739 38112
rect 14803 38048 14819 38112
rect 14883 38048 14899 38112
rect 14963 38048 14969 38112
rect 15840 38088 16000 38118
rect 14653 38047 14969 38048
rect 13813 37906 13879 37909
rect 15840 37906 16000 37936
rect 13813 37904 16000 37906
rect 13813 37848 13818 37904
rect 13874 37848 16000 37904
rect 13813 37846 16000 37848
rect 13813 37843 13879 37846
rect 15840 37816 16000 37846
rect 0 37634 160 37664
rect 749 37634 815 37637
rect 0 37632 815 37634
rect 0 37576 754 37632
rect 810 37576 815 37632
rect 0 37574 815 37576
rect 0 37544 160 37574
rect 749 37571 815 37574
rect 14365 37634 14431 37637
rect 15840 37634 16000 37664
rect 14365 37632 16000 37634
rect 14365 37576 14370 37632
rect 14426 37576 16000 37632
rect 14365 37574 16000 37576
rect 14365 37571 14431 37574
rect 2659 37568 2975 37569
rect 2659 37504 2665 37568
rect 2729 37504 2745 37568
rect 2809 37504 2825 37568
rect 2889 37504 2905 37568
rect 2969 37504 2975 37568
rect 2659 37503 2975 37504
rect 6086 37568 6402 37569
rect 6086 37504 6092 37568
rect 6156 37504 6172 37568
rect 6236 37504 6252 37568
rect 6316 37504 6332 37568
rect 6396 37504 6402 37568
rect 6086 37503 6402 37504
rect 9513 37568 9829 37569
rect 9513 37504 9519 37568
rect 9583 37504 9599 37568
rect 9663 37504 9679 37568
rect 9743 37504 9759 37568
rect 9823 37504 9829 37568
rect 9513 37503 9829 37504
rect 12940 37568 13256 37569
rect 12940 37504 12946 37568
rect 13010 37504 13026 37568
rect 13090 37504 13106 37568
rect 13170 37504 13186 37568
rect 13250 37504 13256 37568
rect 15840 37544 16000 37574
rect 12940 37503 13256 37504
rect 13997 37362 14063 37365
rect 15840 37362 16000 37392
rect 13997 37360 16000 37362
rect 13997 37304 14002 37360
rect 14058 37304 16000 37360
rect 13997 37302 16000 37304
rect 13997 37299 14063 37302
rect 15840 37272 16000 37302
rect 9857 37226 9923 37229
rect 13077 37226 13143 37229
rect 9857 37224 13143 37226
rect 9857 37168 9862 37224
rect 9918 37168 13082 37224
rect 13138 37168 13143 37224
rect 9857 37166 13143 37168
rect 9857 37163 9923 37166
rect 13077 37163 13143 37166
rect 15101 37226 15167 37229
rect 15101 37224 15210 37226
rect 15101 37168 15106 37224
rect 15162 37168 15210 37224
rect 15101 37163 15210 37168
rect 15150 37090 15210 37163
rect 15840 37090 16000 37120
rect 15150 37030 16000 37090
rect 4372 37024 4688 37025
rect 4372 36960 4378 37024
rect 4442 36960 4458 37024
rect 4522 36960 4538 37024
rect 4602 36960 4618 37024
rect 4682 36960 4688 37024
rect 4372 36959 4688 36960
rect 7799 37024 8115 37025
rect 7799 36960 7805 37024
rect 7869 36960 7885 37024
rect 7949 36960 7965 37024
rect 8029 36960 8045 37024
rect 8109 36960 8115 37024
rect 7799 36959 8115 36960
rect 11226 37024 11542 37025
rect 11226 36960 11232 37024
rect 11296 36960 11312 37024
rect 11376 36960 11392 37024
rect 11456 36960 11472 37024
rect 11536 36960 11542 37024
rect 11226 36959 11542 36960
rect 14653 37024 14969 37025
rect 14653 36960 14659 37024
rect 14723 36960 14739 37024
rect 14803 36960 14819 37024
rect 14883 36960 14899 37024
rect 14963 36960 14969 37024
rect 15840 37000 16000 37030
rect 14653 36959 14969 36960
rect 0 36818 160 36848
rect 749 36818 815 36821
rect 0 36816 815 36818
rect 0 36760 754 36816
rect 810 36760 815 36816
rect 0 36758 815 36760
rect 0 36728 160 36758
rect 749 36755 815 36758
rect 13721 36818 13787 36821
rect 15840 36818 16000 36848
rect 13721 36816 16000 36818
rect 13721 36760 13726 36816
rect 13782 36760 16000 36816
rect 13721 36758 16000 36760
rect 13721 36755 13787 36758
rect 15840 36728 16000 36758
rect 6821 36682 6887 36685
rect 13445 36682 13511 36685
rect 6821 36680 13511 36682
rect 6821 36624 6826 36680
rect 6882 36624 13450 36680
rect 13506 36624 13511 36680
rect 6821 36622 13511 36624
rect 6821 36619 6887 36622
rect 13445 36619 13511 36622
rect 14365 36546 14431 36549
rect 15840 36546 16000 36576
rect 14365 36544 16000 36546
rect 14365 36488 14370 36544
rect 14426 36488 16000 36544
rect 14365 36486 16000 36488
rect 14365 36483 14431 36486
rect 2659 36480 2975 36481
rect 2659 36416 2665 36480
rect 2729 36416 2745 36480
rect 2809 36416 2825 36480
rect 2889 36416 2905 36480
rect 2969 36416 2975 36480
rect 2659 36415 2975 36416
rect 6086 36480 6402 36481
rect 6086 36416 6092 36480
rect 6156 36416 6172 36480
rect 6236 36416 6252 36480
rect 6316 36416 6332 36480
rect 6396 36416 6402 36480
rect 6086 36415 6402 36416
rect 9513 36480 9829 36481
rect 9513 36416 9519 36480
rect 9583 36416 9599 36480
rect 9663 36416 9679 36480
rect 9743 36416 9759 36480
rect 9823 36416 9829 36480
rect 9513 36415 9829 36416
rect 12940 36480 13256 36481
rect 12940 36416 12946 36480
rect 13010 36416 13026 36480
rect 13090 36416 13106 36480
rect 13170 36416 13186 36480
rect 13250 36416 13256 36480
rect 15840 36456 16000 36486
rect 12940 36415 13256 36416
rect 10041 36274 10107 36277
rect 13261 36274 13327 36277
rect 10041 36272 13327 36274
rect 10041 36216 10046 36272
rect 10102 36216 13266 36272
rect 13322 36216 13327 36272
rect 10041 36214 13327 36216
rect 10041 36211 10107 36214
rect 13261 36211 13327 36214
rect 13813 36274 13879 36277
rect 15840 36274 16000 36304
rect 13813 36272 16000 36274
rect 13813 36216 13818 36272
rect 13874 36216 16000 36272
rect 13813 36214 16000 36216
rect 13813 36211 13879 36214
rect 15840 36184 16000 36214
rect 10961 36138 11027 36141
rect 13721 36138 13787 36141
rect 10961 36136 13787 36138
rect 10961 36080 10966 36136
rect 11022 36080 13726 36136
rect 13782 36080 13787 36136
rect 10961 36078 13787 36080
rect 10961 36075 11027 36078
rect 13721 36075 13787 36078
rect 0 36002 160 36032
rect 749 36002 815 36005
rect 0 36000 815 36002
rect 0 35944 754 36000
rect 810 35944 815 36000
rect 0 35942 815 35944
rect 0 35912 160 35942
rect 749 35939 815 35942
rect 10501 36004 10567 36005
rect 10501 36000 10548 36004
rect 10612 36002 10618 36004
rect 15101 36002 15167 36005
rect 15840 36002 16000 36032
rect 10501 35944 10506 36000
rect 10501 35940 10548 35944
rect 10612 35942 10658 36002
rect 15101 36000 16000 36002
rect 15101 35944 15106 36000
rect 15162 35944 16000 36000
rect 15101 35942 16000 35944
rect 10612 35940 10618 35942
rect 10501 35939 10567 35940
rect 15101 35939 15167 35942
rect 4372 35936 4688 35937
rect 4372 35872 4378 35936
rect 4442 35872 4458 35936
rect 4522 35872 4538 35936
rect 4602 35872 4618 35936
rect 4682 35872 4688 35936
rect 4372 35871 4688 35872
rect 7799 35936 8115 35937
rect 7799 35872 7805 35936
rect 7869 35872 7885 35936
rect 7949 35872 7965 35936
rect 8029 35872 8045 35936
rect 8109 35872 8115 35936
rect 7799 35871 8115 35872
rect 11226 35936 11542 35937
rect 11226 35872 11232 35936
rect 11296 35872 11312 35936
rect 11376 35872 11392 35936
rect 11456 35872 11472 35936
rect 11536 35872 11542 35936
rect 11226 35871 11542 35872
rect 14653 35936 14969 35937
rect 14653 35872 14659 35936
rect 14723 35872 14739 35936
rect 14803 35872 14819 35936
rect 14883 35872 14899 35936
rect 14963 35872 14969 35936
rect 15840 35912 16000 35942
rect 14653 35871 14969 35872
rect 15377 35866 15443 35869
rect 15377 35864 15578 35866
rect 15377 35808 15382 35864
rect 15438 35808 15578 35864
rect 15377 35806 15578 35808
rect 15377 35803 15443 35806
rect 13261 35730 13327 35733
rect 15518 35730 15578 35806
rect 15840 35730 16000 35760
rect 13261 35728 14474 35730
rect 13261 35672 13266 35728
rect 13322 35672 14474 35728
rect 13261 35670 14474 35672
rect 15518 35670 16000 35730
rect 13261 35667 13327 35670
rect 14414 35458 14474 35670
rect 15840 35640 16000 35670
rect 15840 35458 16000 35488
rect 14414 35398 16000 35458
rect 2659 35392 2975 35393
rect 2659 35328 2665 35392
rect 2729 35328 2745 35392
rect 2809 35328 2825 35392
rect 2889 35328 2905 35392
rect 2969 35328 2975 35392
rect 2659 35327 2975 35328
rect 6086 35392 6402 35393
rect 6086 35328 6092 35392
rect 6156 35328 6172 35392
rect 6236 35328 6252 35392
rect 6316 35328 6332 35392
rect 6396 35328 6402 35392
rect 6086 35327 6402 35328
rect 9513 35392 9829 35393
rect 9513 35328 9519 35392
rect 9583 35328 9599 35392
rect 9663 35328 9679 35392
rect 9743 35328 9759 35392
rect 9823 35328 9829 35392
rect 9513 35327 9829 35328
rect 12940 35392 13256 35393
rect 12940 35328 12946 35392
rect 13010 35328 13026 35392
rect 13090 35328 13106 35392
rect 13170 35328 13186 35392
rect 13250 35328 13256 35392
rect 15840 35368 16000 35398
rect 12940 35327 13256 35328
rect 0 35186 160 35216
rect 749 35186 815 35189
rect 0 35184 815 35186
rect 0 35128 754 35184
rect 810 35128 815 35184
rect 0 35126 815 35128
rect 0 35096 160 35126
rect 749 35123 815 35126
rect 5993 35186 6059 35189
rect 12525 35186 12591 35189
rect 5993 35184 12591 35186
rect 5993 35128 5998 35184
rect 6054 35128 12530 35184
rect 12586 35128 12591 35184
rect 5993 35126 12591 35128
rect 5993 35123 6059 35126
rect 12525 35123 12591 35126
rect 14457 35186 14523 35189
rect 15840 35186 16000 35216
rect 14457 35184 16000 35186
rect 14457 35128 14462 35184
rect 14518 35128 16000 35184
rect 14457 35126 16000 35128
rect 14457 35123 14523 35126
rect 15840 35096 16000 35126
rect 10501 35050 10567 35053
rect 13629 35050 13695 35053
rect 10501 35048 13695 35050
rect 10501 34992 10506 35048
rect 10562 34992 13634 35048
rect 13690 34992 13695 35048
rect 10501 34990 13695 34992
rect 10501 34987 10567 34990
rect 13629 34987 13695 34990
rect 15101 34914 15167 34917
rect 15840 34914 16000 34944
rect 15101 34912 16000 34914
rect 15101 34856 15106 34912
rect 15162 34856 16000 34912
rect 15101 34854 16000 34856
rect 15101 34851 15167 34854
rect 4372 34848 4688 34849
rect 4372 34784 4378 34848
rect 4442 34784 4458 34848
rect 4522 34784 4538 34848
rect 4602 34784 4618 34848
rect 4682 34784 4688 34848
rect 4372 34783 4688 34784
rect 7799 34848 8115 34849
rect 7799 34784 7805 34848
rect 7869 34784 7885 34848
rect 7949 34784 7965 34848
rect 8029 34784 8045 34848
rect 8109 34784 8115 34848
rect 7799 34783 8115 34784
rect 11226 34848 11542 34849
rect 11226 34784 11232 34848
rect 11296 34784 11312 34848
rect 11376 34784 11392 34848
rect 11456 34784 11472 34848
rect 11536 34784 11542 34848
rect 11226 34783 11542 34784
rect 14653 34848 14969 34849
rect 14653 34784 14659 34848
rect 14723 34784 14739 34848
rect 14803 34784 14819 34848
rect 14883 34784 14899 34848
rect 14963 34784 14969 34848
rect 15840 34824 16000 34854
rect 14653 34783 14969 34784
rect 10685 34642 10751 34645
rect 13537 34642 13603 34645
rect 10685 34640 13603 34642
rect 10685 34584 10690 34640
rect 10746 34584 13542 34640
rect 13598 34584 13603 34640
rect 10685 34582 13603 34584
rect 10685 34579 10751 34582
rect 13537 34579 13603 34582
rect 13813 34642 13879 34645
rect 15840 34642 16000 34672
rect 13813 34640 16000 34642
rect 13813 34584 13818 34640
rect 13874 34584 16000 34640
rect 13813 34582 16000 34584
rect 13813 34579 13879 34582
rect 15840 34552 16000 34582
rect 1393 34506 1459 34509
rect 752 34504 1459 34506
rect 752 34448 1398 34504
rect 1454 34448 1459 34504
rect 752 34446 1459 34448
rect 0 34370 160 34400
rect 752 34370 812 34446
rect 1393 34443 1459 34446
rect 12249 34506 12315 34509
rect 15377 34506 15443 34509
rect 12249 34504 15443 34506
rect 12249 34448 12254 34504
rect 12310 34448 15382 34504
rect 15438 34448 15443 34504
rect 12249 34446 15443 34448
rect 12249 34443 12315 34446
rect 15377 34443 15443 34446
rect 15561 34506 15627 34509
rect 15561 34504 15762 34506
rect 15561 34448 15566 34504
rect 15622 34448 15762 34504
rect 15561 34446 15762 34448
rect 15561 34443 15627 34446
rect 0 34310 812 34370
rect 15702 34370 15762 34446
rect 15840 34370 16000 34400
rect 15702 34310 16000 34370
rect 0 34280 160 34310
rect 2659 34304 2975 34305
rect 2659 34240 2665 34304
rect 2729 34240 2745 34304
rect 2809 34240 2825 34304
rect 2889 34240 2905 34304
rect 2969 34240 2975 34304
rect 2659 34239 2975 34240
rect 6086 34304 6402 34305
rect 6086 34240 6092 34304
rect 6156 34240 6172 34304
rect 6236 34240 6252 34304
rect 6316 34240 6332 34304
rect 6396 34240 6402 34304
rect 6086 34239 6402 34240
rect 9513 34304 9829 34305
rect 9513 34240 9519 34304
rect 9583 34240 9599 34304
rect 9663 34240 9679 34304
rect 9743 34240 9759 34304
rect 9823 34240 9829 34304
rect 9513 34239 9829 34240
rect 12940 34304 13256 34305
rect 12940 34240 12946 34304
rect 13010 34240 13026 34304
rect 13090 34240 13106 34304
rect 13170 34240 13186 34304
rect 13250 34240 13256 34304
rect 15840 34280 16000 34310
rect 12940 34239 13256 34240
rect 13261 34098 13327 34101
rect 15840 34098 16000 34128
rect 13261 34096 16000 34098
rect 13261 34040 13266 34096
rect 13322 34040 16000 34096
rect 13261 34038 16000 34040
rect 13261 34035 13327 34038
rect 15840 34008 16000 34038
rect 11513 33962 11579 33965
rect 11646 33962 11652 33964
rect 11513 33960 11652 33962
rect 11513 33904 11518 33960
rect 11574 33904 11652 33960
rect 11513 33902 11652 33904
rect 11513 33899 11579 33902
rect 11646 33900 11652 33902
rect 11716 33900 11722 33964
rect 14549 33962 14615 33965
rect 15377 33962 15443 33965
rect 14549 33960 15210 33962
rect 14549 33904 14554 33960
rect 14610 33904 15210 33960
rect 14549 33902 15210 33904
rect 14549 33899 14615 33902
rect 4372 33760 4688 33761
rect 4372 33696 4378 33760
rect 4442 33696 4458 33760
rect 4522 33696 4538 33760
rect 4602 33696 4618 33760
rect 4682 33696 4688 33760
rect 4372 33695 4688 33696
rect 7799 33760 8115 33761
rect 7799 33696 7805 33760
rect 7869 33696 7885 33760
rect 7949 33696 7965 33760
rect 8029 33696 8045 33760
rect 8109 33696 8115 33760
rect 7799 33695 8115 33696
rect 11226 33760 11542 33761
rect 11226 33696 11232 33760
rect 11296 33696 11312 33760
rect 11376 33696 11392 33760
rect 11456 33696 11472 33760
rect 11536 33696 11542 33760
rect 11226 33695 11542 33696
rect 14653 33760 14969 33761
rect 14653 33696 14659 33760
rect 14723 33696 14739 33760
rect 14803 33696 14819 33760
rect 14883 33696 14899 33760
rect 14963 33696 14969 33760
rect 14653 33695 14969 33696
rect 13486 33628 13492 33692
rect 13556 33690 13562 33692
rect 13629 33690 13695 33693
rect 13556 33688 13695 33690
rect 13556 33632 13634 33688
rect 13690 33632 13695 33688
rect 13556 33630 13695 33632
rect 13556 33628 13562 33630
rect 13629 33627 13695 33630
rect 0 33554 160 33584
rect 749 33554 815 33557
rect 0 33552 815 33554
rect 0 33496 754 33552
rect 810 33496 815 33552
rect 0 33494 815 33496
rect 15150 33554 15210 33902
rect 15377 33960 15578 33962
rect 15377 33904 15382 33960
rect 15438 33904 15578 33960
rect 15377 33902 15578 33904
rect 15377 33899 15443 33902
rect 15518 33826 15578 33902
rect 15840 33826 16000 33856
rect 15518 33766 16000 33826
rect 15840 33736 16000 33766
rect 15840 33554 16000 33584
rect 15150 33494 16000 33554
rect 0 33464 160 33494
rect 749 33491 815 33494
rect 15840 33464 16000 33494
rect 12157 33418 12223 33421
rect 8894 33416 12223 33418
rect 8894 33360 12162 33416
rect 12218 33360 12223 33416
rect 8894 33358 12223 33360
rect 8894 33284 8954 33358
rect 12157 33355 12223 33358
rect 8886 33220 8892 33284
rect 8956 33220 8962 33284
rect 13813 33282 13879 33285
rect 15840 33282 16000 33312
rect 13813 33280 16000 33282
rect 13813 33224 13818 33280
rect 13874 33224 16000 33280
rect 13813 33222 16000 33224
rect 13813 33219 13879 33222
rect 2659 33216 2975 33217
rect 2659 33152 2665 33216
rect 2729 33152 2745 33216
rect 2809 33152 2825 33216
rect 2889 33152 2905 33216
rect 2969 33152 2975 33216
rect 2659 33151 2975 33152
rect 6086 33216 6402 33217
rect 6086 33152 6092 33216
rect 6156 33152 6172 33216
rect 6236 33152 6252 33216
rect 6316 33152 6332 33216
rect 6396 33152 6402 33216
rect 6086 33151 6402 33152
rect 9513 33216 9829 33217
rect 9513 33152 9519 33216
rect 9583 33152 9599 33216
rect 9663 33152 9679 33216
rect 9743 33152 9759 33216
rect 9823 33152 9829 33216
rect 9513 33151 9829 33152
rect 12940 33216 13256 33217
rect 12940 33152 12946 33216
rect 13010 33152 13026 33216
rect 13090 33152 13106 33216
rect 13170 33152 13186 33216
rect 13250 33152 13256 33216
rect 15840 33192 16000 33222
rect 12940 33151 13256 33152
rect 13353 33146 13419 33149
rect 13353 33144 13554 33146
rect 13353 33088 13358 33144
rect 13414 33088 13554 33144
rect 13353 33086 13554 33088
rect 13353 33083 13419 33086
rect 13494 32874 13554 33086
rect 13629 33010 13695 33013
rect 15840 33010 16000 33040
rect 13629 33008 16000 33010
rect 13629 32952 13634 33008
rect 13690 32952 16000 33008
rect 13629 32950 16000 32952
rect 13629 32947 13695 32950
rect 15840 32920 16000 32950
rect 13494 32814 15210 32874
rect 0 32738 160 32768
rect 749 32738 815 32741
rect 0 32736 815 32738
rect 0 32680 754 32736
rect 810 32680 815 32736
rect 0 32678 815 32680
rect 0 32648 160 32678
rect 749 32675 815 32678
rect 12750 32676 12756 32740
rect 12820 32738 12826 32740
rect 14181 32738 14247 32741
rect 12820 32736 14247 32738
rect 12820 32680 14186 32736
rect 14242 32680 14247 32736
rect 12820 32678 14247 32680
rect 15150 32738 15210 32814
rect 15840 32738 16000 32768
rect 15150 32678 16000 32738
rect 12820 32676 12826 32678
rect 14181 32675 14247 32678
rect 4372 32672 4688 32673
rect 4372 32608 4378 32672
rect 4442 32608 4458 32672
rect 4522 32608 4538 32672
rect 4602 32608 4618 32672
rect 4682 32608 4688 32672
rect 4372 32607 4688 32608
rect 7799 32672 8115 32673
rect 7799 32608 7805 32672
rect 7869 32608 7885 32672
rect 7949 32608 7965 32672
rect 8029 32608 8045 32672
rect 8109 32608 8115 32672
rect 7799 32607 8115 32608
rect 11226 32672 11542 32673
rect 11226 32608 11232 32672
rect 11296 32608 11312 32672
rect 11376 32608 11392 32672
rect 11456 32608 11472 32672
rect 11536 32608 11542 32672
rect 11226 32607 11542 32608
rect 14653 32672 14969 32673
rect 14653 32608 14659 32672
rect 14723 32608 14739 32672
rect 14803 32608 14819 32672
rect 14883 32608 14899 32672
rect 14963 32608 14969 32672
rect 15840 32648 16000 32678
rect 14653 32607 14969 32608
rect 12617 32604 12683 32605
rect 12566 32540 12572 32604
rect 12636 32602 12683 32604
rect 12636 32600 12728 32602
rect 12678 32544 12728 32600
rect 12636 32542 12728 32544
rect 12636 32540 12683 32542
rect 12617 32539 12683 32540
rect 12341 32466 12407 32469
rect 15840 32466 16000 32496
rect 12341 32464 16000 32466
rect 12341 32408 12346 32464
rect 12402 32408 16000 32464
rect 12341 32406 16000 32408
rect 12341 32403 12407 32406
rect 15840 32376 16000 32406
rect 6913 32330 6979 32333
rect 12985 32330 13051 32333
rect 6913 32328 13051 32330
rect 6913 32272 6918 32328
rect 6974 32272 12990 32328
rect 13046 32272 13051 32328
rect 6913 32270 13051 32272
rect 6913 32267 6979 32270
rect 12985 32267 13051 32270
rect 13997 32330 14063 32333
rect 13997 32328 14290 32330
rect 13997 32272 14002 32328
rect 14058 32272 14290 32328
rect 13997 32270 14290 32272
rect 13997 32267 14063 32270
rect 2659 32128 2975 32129
rect 2659 32064 2665 32128
rect 2729 32064 2745 32128
rect 2809 32064 2825 32128
rect 2889 32064 2905 32128
rect 2969 32064 2975 32128
rect 2659 32063 2975 32064
rect 6086 32128 6402 32129
rect 6086 32064 6092 32128
rect 6156 32064 6172 32128
rect 6236 32064 6252 32128
rect 6316 32064 6332 32128
rect 6396 32064 6402 32128
rect 6086 32063 6402 32064
rect 9513 32128 9829 32129
rect 9513 32064 9519 32128
rect 9583 32064 9599 32128
rect 9663 32064 9679 32128
rect 9743 32064 9759 32128
rect 9823 32064 9829 32128
rect 9513 32063 9829 32064
rect 12940 32128 13256 32129
rect 12940 32064 12946 32128
rect 13010 32064 13026 32128
rect 13090 32064 13106 32128
rect 13170 32064 13186 32128
rect 13250 32064 13256 32128
rect 12940 32063 13256 32064
rect 0 31922 160 31952
rect 749 31922 815 31925
rect 0 31920 815 31922
rect 0 31864 754 31920
rect 810 31864 815 31920
rect 0 31862 815 31864
rect 0 31832 160 31862
rect 749 31859 815 31862
rect 7230 31860 7236 31924
rect 7300 31922 7306 31924
rect 11053 31922 11119 31925
rect 7300 31920 11119 31922
rect 7300 31864 11058 31920
rect 11114 31864 11119 31920
rect 7300 31862 11119 31864
rect 7300 31860 7306 31862
rect 11053 31859 11119 31862
rect 11513 31922 11579 31925
rect 13813 31922 13879 31925
rect 11513 31920 13879 31922
rect 11513 31864 11518 31920
rect 11574 31864 13818 31920
rect 13874 31864 13879 31920
rect 11513 31862 13879 31864
rect 14230 31922 14290 32270
rect 15561 32194 15627 32197
rect 15840 32194 16000 32224
rect 15561 32192 16000 32194
rect 15561 32136 15566 32192
rect 15622 32136 16000 32192
rect 15561 32134 16000 32136
rect 15561 32131 15627 32134
rect 15840 32104 16000 32134
rect 15840 31922 16000 31952
rect 14230 31862 16000 31922
rect 11513 31859 11579 31862
rect 13813 31859 13879 31862
rect 15840 31832 16000 31862
rect 11973 31786 12039 31789
rect 14038 31786 14044 31788
rect 11973 31784 14044 31786
rect 11973 31728 11978 31784
rect 12034 31728 14044 31784
rect 11973 31726 14044 31728
rect 11973 31723 12039 31726
rect 14038 31724 14044 31726
rect 14108 31724 14114 31788
rect 15469 31650 15535 31653
rect 15840 31650 16000 31680
rect 15469 31648 16000 31650
rect 15469 31592 15474 31648
rect 15530 31592 16000 31648
rect 15469 31590 16000 31592
rect 15469 31587 15535 31590
rect 4372 31584 4688 31585
rect 4372 31520 4378 31584
rect 4442 31520 4458 31584
rect 4522 31520 4538 31584
rect 4602 31520 4618 31584
rect 4682 31520 4688 31584
rect 4372 31519 4688 31520
rect 7799 31584 8115 31585
rect 7799 31520 7805 31584
rect 7869 31520 7885 31584
rect 7949 31520 7965 31584
rect 8029 31520 8045 31584
rect 8109 31520 8115 31584
rect 7799 31519 8115 31520
rect 11226 31584 11542 31585
rect 11226 31520 11232 31584
rect 11296 31520 11312 31584
rect 11376 31520 11392 31584
rect 11456 31520 11472 31584
rect 11536 31520 11542 31584
rect 11226 31519 11542 31520
rect 14653 31584 14969 31585
rect 14653 31520 14659 31584
rect 14723 31520 14739 31584
rect 14803 31520 14819 31584
rect 14883 31520 14899 31584
rect 14963 31520 14969 31584
rect 15840 31560 16000 31590
rect 14653 31519 14969 31520
rect 11881 31378 11947 31381
rect 12341 31378 12407 31381
rect 15840 31378 16000 31408
rect 11881 31376 12407 31378
rect 11881 31320 11886 31376
rect 11942 31320 12346 31376
rect 12402 31320 12407 31376
rect 11881 31318 12407 31320
rect 11881 31315 11947 31318
rect 12341 31315 12407 31318
rect 15564 31318 16000 31378
rect 13353 31242 13419 31245
rect 15564 31242 15624 31318
rect 15840 31288 16000 31318
rect 13353 31240 15624 31242
rect 13353 31184 13358 31240
rect 13414 31184 15624 31240
rect 13353 31182 15624 31184
rect 13353 31179 13419 31182
rect 0 31106 160 31136
rect 749 31106 815 31109
rect 15840 31106 16000 31136
rect 0 31104 815 31106
rect 0 31048 754 31104
rect 810 31048 815 31104
rect 0 31046 815 31048
rect 0 31016 160 31046
rect 749 31043 815 31046
rect 14230 31046 16000 31106
rect 2659 31040 2975 31041
rect 2659 30976 2665 31040
rect 2729 30976 2745 31040
rect 2809 30976 2825 31040
rect 2889 30976 2905 31040
rect 2969 30976 2975 31040
rect 2659 30975 2975 30976
rect 6086 31040 6402 31041
rect 6086 30976 6092 31040
rect 6156 30976 6172 31040
rect 6236 30976 6252 31040
rect 6316 30976 6332 31040
rect 6396 30976 6402 31040
rect 6086 30975 6402 30976
rect 9513 31040 9829 31041
rect 9513 30976 9519 31040
rect 9583 30976 9599 31040
rect 9663 30976 9679 31040
rect 9743 30976 9759 31040
rect 9823 30976 9829 31040
rect 9513 30975 9829 30976
rect 12940 31040 13256 31041
rect 12940 30976 12946 31040
rect 13010 30976 13026 31040
rect 13090 30976 13106 31040
rect 13170 30976 13186 31040
rect 13250 30976 13256 31040
rect 12940 30975 13256 30976
rect 9070 30772 9076 30836
rect 9140 30834 9146 30836
rect 11237 30834 11303 30837
rect 9140 30832 11303 30834
rect 9140 30776 11242 30832
rect 11298 30776 11303 30832
rect 9140 30774 11303 30776
rect 9140 30772 9146 30774
rect 11237 30771 11303 30774
rect 12157 30834 12223 30837
rect 14230 30834 14290 31046
rect 15840 31016 16000 31046
rect 12157 30832 14290 30834
rect 12157 30776 12162 30832
rect 12218 30776 14290 30832
rect 12157 30774 14290 30776
rect 14549 30834 14615 30837
rect 15840 30834 16000 30864
rect 14549 30832 16000 30834
rect 14549 30776 14554 30832
rect 14610 30776 16000 30832
rect 14549 30774 16000 30776
rect 12157 30771 12223 30774
rect 14549 30771 14615 30774
rect 15840 30744 16000 30774
rect 10726 30636 10732 30700
rect 10796 30698 10802 30700
rect 14273 30698 14339 30701
rect 10796 30696 14339 30698
rect 10796 30640 14278 30696
rect 14334 30640 14339 30696
rect 10796 30638 14339 30640
rect 10796 30636 10802 30638
rect 14273 30635 14339 30638
rect 13537 30562 13603 30565
rect 15653 30562 15719 30565
rect 15840 30562 16000 30592
rect 13537 30560 14428 30562
rect 13537 30504 13542 30560
rect 13598 30504 14428 30560
rect 13537 30502 14428 30504
rect 13537 30499 13603 30502
rect 4372 30496 4688 30497
rect 4372 30432 4378 30496
rect 4442 30432 4458 30496
rect 4522 30432 4538 30496
rect 4602 30432 4618 30496
rect 4682 30432 4688 30496
rect 4372 30431 4688 30432
rect 7799 30496 8115 30497
rect 7799 30432 7805 30496
rect 7869 30432 7885 30496
rect 7949 30432 7965 30496
rect 8029 30432 8045 30496
rect 8109 30432 8115 30496
rect 7799 30431 8115 30432
rect 11226 30496 11542 30497
rect 11226 30432 11232 30496
rect 11296 30432 11312 30496
rect 11376 30432 11392 30496
rect 11456 30432 11472 30496
rect 11536 30432 11542 30496
rect 11226 30431 11542 30432
rect 0 30290 160 30320
rect 1393 30290 1459 30293
rect 0 30288 1459 30290
rect 0 30232 1398 30288
rect 1454 30232 1459 30288
rect 0 30230 1459 30232
rect 0 30200 160 30230
rect 1393 30227 1459 30230
rect 11605 30290 11671 30293
rect 14368 30290 14428 30502
rect 15653 30560 16000 30562
rect 15653 30504 15658 30560
rect 15714 30504 16000 30560
rect 15653 30502 16000 30504
rect 15653 30499 15719 30502
rect 14653 30496 14969 30497
rect 14653 30432 14659 30496
rect 14723 30432 14739 30496
rect 14803 30432 14819 30496
rect 14883 30432 14899 30496
rect 14963 30432 14969 30496
rect 15840 30472 16000 30502
rect 14653 30431 14969 30432
rect 15840 30290 16000 30320
rect 11605 30288 14244 30290
rect 11605 30232 11610 30288
rect 11666 30232 14244 30288
rect 11605 30230 14244 30232
rect 14368 30230 16000 30290
rect 11605 30227 11671 30230
rect 12249 30154 12315 30157
rect 12566 30154 12572 30156
rect 12249 30152 12572 30154
rect 12249 30096 12254 30152
rect 12310 30096 12572 30152
rect 12249 30094 12572 30096
rect 12249 30091 12315 30094
rect 12566 30092 12572 30094
rect 12636 30092 12642 30156
rect 12758 30094 14106 30154
rect 10777 30018 10843 30021
rect 11145 30018 11211 30021
rect 10777 30016 11211 30018
rect 10777 29960 10782 30016
rect 10838 29960 11150 30016
rect 11206 29960 11211 30016
rect 10777 29958 11211 29960
rect 10777 29955 10843 29958
rect 11145 29955 11211 29958
rect 11329 30018 11395 30021
rect 12758 30018 12818 30094
rect 11329 30016 12818 30018
rect 11329 29960 11334 30016
rect 11390 29960 12818 30016
rect 11329 29958 12818 29960
rect 11329 29955 11395 29958
rect 2659 29952 2975 29953
rect 2659 29888 2665 29952
rect 2729 29888 2745 29952
rect 2809 29888 2825 29952
rect 2889 29888 2905 29952
rect 2969 29888 2975 29952
rect 2659 29887 2975 29888
rect 6086 29952 6402 29953
rect 6086 29888 6092 29952
rect 6156 29888 6172 29952
rect 6236 29888 6252 29952
rect 6316 29888 6332 29952
rect 6396 29888 6402 29952
rect 6086 29887 6402 29888
rect 9513 29952 9829 29953
rect 9513 29888 9519 29952
rect 9583 29888 9599 29952
rect 9663 29888 9679 29952
rect 9743 29888 9759 29952
rect 9823 29888 9829 29952
rect 9513 29887 9829 29888
rect 12940 29952 13256 29953
rect 12940 29888 12946 29952
rect 13010 29888 13026 29952
rect 13090 29888 13106 29952
rect 13170 29888 13186 29952
rect 13250 29888 13256 29952
rect 12940 29887 13256 29888
rect 10685 29882 10751 29885
rect 11421 29882 11487 29885
rect 10685 29880 11487 29882
rect 10685 29824 10690 29880
rect 10746 29824 11426 29880
rect 11482 29824 11487 29880
rect 10685 29822 11487 29824
rect 10685 29819 10751 29822
rect 11421 29819 11487 29822
rect 12341 29882 12407 29885
rect 12750 29882 12756 29884
rect 12341 29880 12756 29882
rect 12341 29824 12346 29880
rect 12402 29824 12756 29880
rect 12341 29822 12756 29824
rect 12341 29819 12407 29822
rect 12750 29820 12756 29822
rect 12820 29820 12826 29884
rect 14046 29882 14106 30094
rect 14184 30018 14244 30230
rect 15840 30200 16000 30230
rect 15840 30018 16000 30048
rect 14184 29958 16000 30018
rect 15840 29928 16000 29958
rect 14046 29822 15394 29882
rect 8569 29746 8635 29749
rect 9581 29746 9647 29749
rect 11237 29746 11303 29749
rect 8569 29744 11303 29746
rect 8569 29688 8574 29744
rect 8630 29688 9586 29744
rect 9642 29688 11242 29744
rect 11298 29688 11303 29744
rect 8569 29686 11303 29688
rect 8569 29683 8635 29686
rect 9581 29683 9647 29686
rect 11237 29683 11303 29686
rect 11789 29746 11855 29749
rect 15334 29746 15394 29822
rect 15840 29746 16000 29776
rect 11789 29744 15210 29746
rect 11789 29688 11794 29744
rect 11850 29688 15210 29744
rect 11789 29686 15210 29688
rect 15334 29686 16000 29746
rect 11789 29683 11855 29686
rect 10726 29548 10732 29612
rect 10796 29610 10802 29612
rect 11237 29610 11303 29613
rect 10796 29608 11303 29610
rect 10796 29552 11242 29608
rect 11298 29552 11303 29608
rect 10796 29550 11303 29552
rect 10796 29548 10802 29550
rect 11237 29547 11303 29550
rect 12617 29608 12683 29613
rect 12617 29552 12622 29608
rect 12678 29552 12683 29608
rect 12617 29547 12683 29552
rect 0 29474 160 29504
rect 749 29474 815 29477
rect 0 29472 815 29474
rect 0 29416 754 29472
rect 810 29416 815 29472
rect 0 29414 815 29416
rect 0 29384 160 29414
rect 749 29411 815 29414
rect 4372 29408 4688 29409
rect 4372 29344 4378 29408
rect 4442 29344 4458 29408
rect 4522 29344 4538 29408
rect 4602 29344 4618 29408
rect 4682 29344 4688 29408
rect 4372 29343 4688 29344
rect 7799 29408 8115 29409
rect 7799 29344 7805 29408
rect 7869 29344 7885 29408
rect 7949 29344 7965 29408
rect 8029 29344 8045 29408
rect 8109 29344 8115 29408
rect 7799 29343 8115 29344
rect 11226 29408 11542 29409
rect 11226 29344 11232 29408
rect 11296 29344 11312 29408
rect 11376 29344 11392 29408
rect 11456 29344 11472 29408
rect 11536 29344 11542 29408
rect 11226 29343 11542 29344
rect 8201 29338 8267 29341
rect 9213 29338 9279 29341
rect 12620 29338 12680 29547
rect 15150 29474 15210 29686
rect 15840 29656 16000 29686
rect 15840 29474 16000 29504
rect 15150 29414 16000 29474
rect 14653 29408 14969 29409
rect 14653 29344 14659 29408
rect 14723 29344 14739 29408
rect 14803 29344 14819 29408
rect 14883 29344 14899 29408
rect 14963 29344 14969 29408
rect 15840 29384 16000 29414
rect 14653 29343 14969 29344
rect 8201 29336 9279 29338
rect 8201 29280 8206 29336
rect 8262 29280 9218 29336
rect 9274 29280 9279 29336
rect 8201 29278 9279 29280
rect 8201 29275 8267 29278
rect 9213 29275 9279 29278
rect 11976 29278 12680 29338
rect 5625 29202 5691 29205
rect 11976 29202 12036 29278
rect 5625 29200 12036 29202
rect 5625 29144 5630 29200
rect 5686 29144 12036 29200
rect 5625 29142 12036 29144
rect 12249 29202 12315 29205
rect 13486 29202 13492 29204
rect 12249 29200 13492 29202
rect 12249 29144 12254 29200
rect 12310 29144 13492 29200
rect 12249 29142 13492 29144
rect 5625 29139 5691 29142
rect 12249 29139 12315 29142
rect 13486 29140 13492 29142
rect 13556 29140 13562 29204
rect 13813 29202 13879 29205
rect 15840 29202 16000 29232
rect 13813 29200 16000 29202
rect 13813 29144 13818 29200
rect 13874 29144 16000 29200
rect 13813 29142 16000 29144
rect 13813 29139 13879 29142
rect 15840 29112 16000 29142
rect 11605 29068 11671 29069
rect 11605 29064 11652 29068
rect 11716 29066 11722 29068
rect 12617 29066 12683 29069
rect 13169 29066 13235 29069
rect 11605 29008 11610 29064
rect 11605 29004 11652 29008
rect 11716 29006 11762 29066
rect 12617 29064 13235 29066
rect 12617 29008 12622 29064
rect 12678 29008 13174 29064
rect 13230 29008 13235 29064
rect 12617 29006 13235 29008
rect 11716 29004 11722 29006
rect 11605 29003 11671 29004
rect 12617 29003 12683 29006
rect 13169 29003 13235 29006
rect 1393 28930 1459 28933
rect 15840 28930 16000 28960
rect 752 28928 1459 28930
rect 752 28872 1398 28928
rect 1454 28872 1459 28928
rect 752 28870 1459 28872
rect 0 28658 160 28688
rect 752 28658 812 28870
rect 1393 28867 1459 28870
rect 14046 28870 16000 28930
rect 2659 28864 2975 28865
rect 2659 28800 2665 28864
rect 2729 28800 2745 28864
rect 2809 28800 2825 28864
rect 2889 28800 2905 28864
rect 2969 28800 2975 28864
rect 2659 28799 2975 28800
rect 6086 28864 6402 28865
rect 6086 28800 6092 28864
rect 6156 28800 6172 28864
rect 6236 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6402 28864
rect 6086 28799 6402 28800
rect 9513 28864 9829 28865
rect 9513 28800 9519 28864
rect 9583 28800 9599 28864
rect 9663 28800 9679 28864
rect 9743 28800 9759 28864
rect 9823 28800 9829 28864
rect 9513 28799 9829 28800
rect 12940 28864 13256 28865
rect 12940 28800 12946 28864
rect 13010 28800 13026 28864
rect 13090 28800 13106 28864
rect 13170 28800 13186 28864
rect 13250 28800 13256 28864
rect 12940 28799 13256 28800
rect 11053 28794 11119 28797
rect 12750 28794 12756 28796
rect 11053 28792 12756 28794
rect 11053 28736 11058 28792
rect 11114 28736 12756 28792
rect 11053 28734 12756 28736
rect 11053 28731 11119 28734
rect 12750 28732 12756 28734
rect 12820 28732 12826 28796
rect 14046 28658 14106 28870
rect 15840 28840 16000 28870
rect 0 28598 812 28658
rect 12390 28598 14106 28658
rect 14273 28658 14339 28661
rect 15840 28658 16000 28688
rect 14273 28656 16000 28658
rect 14273 28600 14278 28656
rect 14334 28600 16000 28656
rect 14273 28598 16000 28600
rect 0 28568 160 28598
rect 1710 28460 1716 28524
rect 1780 28522 1786 28524
rect 9213 28522 9279 28525
rect 1780 28520 9279 28522
rect 1780 28464 9218 28520
rect 9274 28464 9279 28520
rect 1780 28462 9279 28464
rect 1780 28460 1786 28462
rect 9213 28459 9279 28462
rect 11053 28522 11119 28525
rect 12390 28522 12450 28598
rect 14273 28595 14339 28598
rect 15840 28568 16000 28598
rect 11053 28520 12450 28522
rect 11053 28464 11058 28520
rect 11114 28464 12450 28520
rect 11053 28462 12450 28464
rect 11053 28459 11119 28462
rect 12750 28460 12756 28524
rect 12820 28522 12826 28524
rect 13813 28522 13879 28525
rect 12820 28520 13879 28522
rect 12820 28464 13818 28520
rect 13874 28464 13879 28520
rect 12820 28462 13879 28464
rect 12820 28460 12826 28462
rect 13813 28459 13879 28462
rect 15561 28386 15627 28389
rect 15840 28386 16000 28416
rect 15561 28384 16000 28386
rect 15561 28328 15566 28384
rect 15622 28328 16000 28384
rect 15561 28326 16000 28328
rect 15561 28323 15627 28326
rect 4372 28320 4688 28321
rect 4372 28256 4378 28320
rect 4442 28256 4458 28320
rect 4522 28256 4538 28320
rect 4602 28256 4618 28320
rect 4682 28256 4688 28320
rect 4372 28255 4688 28256
rect 7799 28320 8115 28321
rect 7799 28256 7805 28320
rect 7869 28256 7885 28320
rect 7949 28256 7965 28320
rect 8029 28256 8045 28320
rect 8109 28256 8115 28320
rect 7799 28255 8115 28256
rect 11226 28320 11542 28321
rect 11226 28256 11232 28320
rect 11296 28256 11312 28320
rect 11376 28256 11392 28320
rect 11456 28256 11472 28320
rect 11536 28256 11542 28320
rect 11226 28255 11542 28256
rect 14653 28320 14969 28321
rect 14653 28256 14659 28320
rect 14723 28256 14739 28320
rect 14803 28256 14819 28320
rect 14883 28256 14899 28320
rect 14963 28256 14969 28320
rect 15840 28296 16000 28326
rect 14653 28255 14969 28256
rect 13854 28250 13860 28252
rect 11654 28190 13860 28250
rect 9581 28114 9647 28117
rect 11654 28114 11714 28190
rect 13854 28188 13860 28190
rect 13924 28188 13930 28252
rect 9581 28112 11714 28114
rect 9581 28056 9586 28112
rect 9642 28056 11714 28112
rect 9581 28054 11714 28056
rect 12341 28114 12407 28117
rect 15840 28114 16000 28144
rect 12341 28112 13554 28114
rect 12341 28056 12346 28112
rect 12402 28056 13554 28112
rect 12341 28054 13554 28056
rect 9581 28051 9647 28054
rect 12341 28051 12407 28054
rect 0 27842 160 27872
rect 749 27842 815 27845
rect 0 27840 815 27842
rect 0 27784 754 27840
rect 810 27784 815 27840
rect 0 27782 815 27784
rect 13494 27842 13554 28054
rect 15702 28054 16000 28114
rect 13629 27978 13695 27981
rect 15702 27978 15762 28054
rect 15840 28024 16000 28054
rect 13629 27976 15762 27978
rect 13629 27920 13634 27976
rect 13690 27920 15762 27976
rect 13629 27918 15762 27920
rect 13629 27915 13695 27918
rect 15840 27842 16000 27872
rect 13494 27782 16000 27842
rect 0 27752 160 27782
rect 749 27779 815 27782
rect 2659 27776 2975 27777
rect 2659 27712 2665 27776
rect 2729 27712 2745 27776
rect 2809 27712 2825 27776
rect 2889 27712 2905 27776
rect 2969 27712 2975 27776
rect 2659 27711 2975 27712
rect 6086 27776 6402 27777
rect 6086 27712 6092 27776
rect 6156 27712 6172 27776
rect 6236 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6402 27776
rect 6086 27711 6402 27712
rect 9513 27776 9829 27777
rect 9513 27712 9519 27776
rect 9583 27712 9599 27776
rect 9663 27712 9679 27776
rect 9743 27712 9759 27776
rect 9823 27712 9829 27776
rect 9513 27711 9829 27712
rect 12940 27776 13256 27777
rect 12940 27712 12946 27776
rect 13010 27712 13026 27776
rect 13090 27712 13106 27776
rect 13170 27712 13186 27776
rect 13250 27712 13256 27776
rect 15840 27752 16000 27782
rect 12940 27711 13256 27712
rect 11973 27570 12039 27573
rect 15469 27570 15535 27573
rect 15840 27570 16000 27600
rect 11973 27568 15210 27570
rect 11973 27512 11978 27568
rect 12034 27512 15210 27568
rect 11973 27510 15210 27512
rect 11973 27507 12039 27510
rect 9857 27434 9923 27437
rect 11513 27434 11579 27437
rect 12433 27434 12499 27437
rect 12709 27434 12775 27437
rect 9857 27432 12775 27434
rect 9857 27376 9862 27432
rect 9918 27376 11518 27432
rect 11574 27376 12438 27432
rect 12494 27376 12714 27432
rect 12770 27376 12775 27432
rect 9857 27374 12775 27376
rect 9857 27371 9923 27374
rect 11513 27371 11579 27374
rect 12433 27371 12499 27374
rect 12709 27371 12775 27374
rect 13670 27372 13676 27436
rect 13740 27434 13746 27436
rect 13813 27434 13879 27437
rect 13740 27432 13879 27434
rect 13740 27376 13818 27432
rect 13874 27376 13879 27432
rect 13740 27374 13879 27376
rect 13740 27372 13746 27374
rect 13813 27371 13879 27374
rect 15150 27298 15210 27510
rect 15469 27568 16000 27570
rect 15469 27512 15474 27568
rect 15530 27512 16000 27568
rect 15469 27510 16000 27512
rect 15469 27507 15535 27510
rect 15840 27480 16000 27510
rect 15840 27298 16000 27328
rect 15150 27238 16000 27298
rect 4372 27232 4688 27233
rect 4372 27168 4378 27232
rect 4442 27168 4458 27232
rect 4522 27168 4538 27232
rect 4602 27168 4618 27232
rect 4682 27168 4688 27232
rect 4372 27167 4688 27168
rect 7799 27232 8115 27233
rect 7799 27168 7805 27232
rect 7869 27168 7885 27232
rect 7949 27168 7965 27232
rect 8029 27168 8045 27232
rect 8109 27168 8115 27232
rect 7799 27167 8115 27168
rect 11226 27232 11542 27233
rect 11226 27168 11232 27232
rect 11296 27168 11312 27232
rect 11376 27168 11392 27232
rect 11456 27168 11472 27232
rect 11536 27168 11542 27232
rect 11226 27167 11542 27168
rect 14653 27232 14969 27233
rect 14653 27168 14659 27232
rect 14723 27168 14739 27232
rect 14803 27168 14819 27232
rect 14883 27168 14899 27232
rect 14963 27168 14969 27232
rect 15840 27208 16000 27238
rect 14653 27167 14969 27168
rect 0 27026 160 27056
rect 749 27026 815 27029
rect 0 27024 815 27026
rect 0 26968 754 27024
rect 810 26968 815 27024
rect 0 26966 815 26968
rect 0 26936 160 26966
rect 749 26963 815 26966
rect 14181 27026 14247 27029
rect 15840 27026 16000 27056
rect 14181 27024 16000 27026
rect 14181 26968 14186 27024
rect 14242 26968 16000 27024
rect 14181 26966 16000 26968
rect 14181 26963 14247 26966
rect 15840 26936 16000 26966
rect 14641 26754 14707 26757
rect 15840 26754 16000 26784
rect 14641 26752 16000 26754
rect 14641 26696 14646 26752
rect 14702 26696 16000 26752
rect 14641 26694 16000 26696
rect 14641 26691 14707 26694
rect 2659 26688 2975 26689
rect 2659 26624 2665 26688
rect 2729 26624 2745 26688
rect 2809 26624 2825 26688
rect 2889 26624 2905 26688
rect 2969 26624 2975 26688
rect 2659 26623 2975 26624
rect 6086 26688 6402 26689
rect 6086 26624 6092 26688
rect 6156 26624 6172 26688
rect 6236 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6402 26688
rect 6086 26623 6402 26624
rect 9513 26688 9829 26689
rect 9513 26624 9519 26688
rect 9583 26624 9599 26688
rect 9663 26624 9679 26688
rect 9743 26624 9759 26688
rect 9823 26624 9829 26688
rect 9513 26623 9829 26624
rect 12940 26688 13256 26689
rect 12940 26624 12946 26688
rect 13010 26624 13026 26688
rect 13090 26624 13106 26688
rect 13170 26624 13186 26688
rect 13250 26624 13256 26688
rect 15840 26664 16000 26694
rect 12940 26623 13256 26624
rect 11881 26482 11947 26485
rect 15840 26482 16000 26512
rect 11881 26480 16000 26482
rect 11881 26424 11886 26480
rect 11942 26424 16000 26480
rect 11881 26422 16000 26424
rect 11881 26419 11947 26422
rect 15840 26392 16000 26422
rect 3918 26284 3924 26348
rect 3988 26346 3994 26348
rect 10133 26346 10199 26349
rect 3988 26344 10199 26346
rect 3988 26288 10138 26344
rect 10194 26288 10199 26344
rect 3988 26286 10199 26288
rect 3988 26284 3994 26286
rect 10133 26283 10199 26286
rect 0 26210 160 26240
rect 1485 26210 1551 26213
rect 0 26208 1551 26210
rect 0 26152 1490 26208
rect 1546 26152 1551 26208
rect 0 26150 1551 26152
rect 0 26120 160 26150
rect 1485 26147 1551 26150
rect 15101 26210 15167 26213
rect 15840 26210 16000 26240
rect 15101 26208 16000 26210
rect 15101 26152 15106 26208
rect 15162 26152 16000 26208
rect 15101 26150 16000 26152
rect 15101 26147 15167 26150
rect 4372 26144 4688 26145
rect 4372 26080 4378 26144
rect 4442 26080 4458 26144
rect 4522 26080 4538 26144
rect 4602 26080 4618 26144
rect 4682 26080 4688 26144
rect 4372 26079 4688 26080
rect 7799 26144 8115 26145
rect 7799 26080 7805 26144
rect 7869 26080 7885 26144
rect 7949 26080 7965 26144
rect 8029 26080 8045 26144
rect 8109 26080 8115 26144
rect 7799 26079 8115 26080
rect 11226 26144 11542 26145
rect 11226 26080 11232 26144
rect 11296 26080 11312 26144
rect 11376 26080 11392 26144
rect 11456 26080 11472 26144
rect 11536 26080 11542 26144
rect 11226 26079 11542 26080
rect 14653 26144 14969 26145
rect 14653 26080 14659 26144
rect 14723 26080 14739 26144
rect 14803 26080 14819 26144
rect 14883 26080 14899 26144
rect 14963 26080 14969 26144
rect 15840 26120 16000 26150
rect 14653 26079 14969 26080
rect 15469 25938 15535 25941
rect 15840 25938 16000 25968
rect 15469 25936 16000 25938
rect 15469 25880 15474 25936
rect 15530 25880 16000 25936
rect 15469 25878 16000 25880
rect 15469 25875 15535 25878
rect 15840 25848 16000 25878
rect 12249 25802 12315 25805
rect 13629 25802 13695 25805
rect 12249 25800 13695 25802
rect 12249 25744 12254 25800
rect 12310 25744 13634 25800
rect 13690 25744 13695 25800
rect 12249 25742 13695 25744
rect 12249 25739 12315 25742
rect 13629 25739 13695 25742
rect 14181 25666 14247 25669
rect 15840 25666 16000 25696
rect 14181 25664 16000 25666
rect 14181 25608 14186 25664
rect 14242 25608 16000 25664
rect 14181 25606 16000 25608
rect 14181 25603 14247 25606
rect 2659 25600 2975 25601
rect 2659 25536 2665 25600
rect 2729 25536 2745 25600
rect 2809 25536 2825 25600
rect 2889 25536 2905 25600
rect 2969 25536 2975 25600
rect 2659 25535 2975 25536
rect 6086 25600 6402 25601
rect 6086 25536 6092 25600
rect 6156 25536 6172 25600
rect 6236 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6402 25600
rect 6086 25535 6402 25536
rect 9513 25600 9829 25601
rect 9513 25536 9519 25600
rect 9583 25536 9599 25600
rect 9663 25536 9679 25600
rect 9743 25536 9759 25600
rect 9823 25536 9829 25600
rect 9513 25535 9829 25536
rect 12940 25600 13256 25601
rect 12940 25536 12946 25600
rect 13010 25536 13026 25600
rect 13090 25536 13106 25600
rect 13170 25536 13186 25600
rect 13250 25536 13256 25600
rect 15840 25576 16000 25606
rect 12940 25535 13256 25536
rect 14549 25530 14615 25533
rect 14549 25528 15762 25530
rect 14549 25472 14554 25528
rect 14610 25472 15762 25528
rect 14549 25470 15762 25472
rect 14549 25467 14615 25470
rect 0 25394 160 25424
rect 749 25394 815 25397
rect 0 25392 815 25394
rect 0 25336 754 25392
rect 810 25336 815 25392
rect 0 25334 815 25336
rect 15702 25394 15762 25470
rect 15840 25394 16000 25424
rect 15702 25334 16000 25394
rect 0 25304 160 25334
rect 749 25331 815 25334
rect 15840 25304 16000 25334
rect 6494 25196 6500 25260
rect 6564 25258 6570 25260
rect 8201 25258 8267 25261
rect 11145 25258 11211 25261
rect 6564 25256 8402 25258
rect 6564 25200 8206 25256
rect 8262 25200 8402 25256
rect 6564 25198 8402 25200
rect 6564 25196 6570 25198
rect 8201 25195 8267 25198
rect 8342 25122 8402 25198
rect 11145 25256 15210 25258
rect 11145 25200 11150 25256
rect 11206 25200 15210 25256
rect 11145 25198 15210 25200
rect 11145 25195 11211 25198
rect 10409 25122 10475 25125
rect 10542 25122 10548 25124
rect 8342 25120 10548 25122
rect 8342 25064 10414 25120
rect 10470 25064 10548 25120
rect 8342 25062 10548 25064
rect 10409 25059 10475 25062
rect 10542 25060 10548 25062
rect 10612 25060 10618 25124
rect 15150 25122 15210 25198
rect 15840 25122 16000 25152
rect 15150 25062 16000 25122
rect 4372 25056 4688 25057
rect 4372 24992 4378 25056
rect 4442 24992 4458 25056
rect 4522 24992 4538 25056
rect 4602 24992 4618 25056
rect 4682 24992 4688 25056
rect 4372 24991 4688 24992
rect 7799 25056 8115 25057
rect 7799 24992 7805 25056
rect 7869 24992 7885 25056
rect 7949 24992 7965 25056
rect 8029 24992 8045 25056
rect 8109 24992 8115 25056
rect 7799 24991 8115 24992
rect 11226 25056 11542 25057
rect 11226 24992 11232 25056
rect 11296 24992 11312 25056
rect 11376 24992 11392 25056
rect 11456 24992 11472 25056
rect 11536 24992 11542 25056
rect 11226 24991 11542 24992
rect 14653 25056 14969 25057
rect 14653 24992 14659 25056
rect 14723 24992 14739 25056
rect 14803 24992 14819 25056
rect 14883 24992 14899 25056
rect 14963 24992 14969 25056
rect 15840 25032 16000 25062
rect 14653 24991 14969 24992
rect 11881 24850 11947 24853
rect 15840 24850 16000 24880
rect 11881 24848 16000 24850
rect 11881 24792 11886 24848
rect 11942 24792 16000 24848
rect 11881 24790 16000 24792
rect 11881 24787 11947 24790
rect 15840 24760 16000 24790
rect 10542 24652 10548 24716
rect 10612 24714 10618 24716
rect 13169 24714 13235 24717
rect 13486 24714 13492 24716
rect 10612 24712 13492 24714
rect 10612 24656 13174 24712
rect 13230 24656 13492 24712
rect 10612 24654 13492 24656
rect 10612 24652 10618 24654
rect 13169 24651 13235 24654
rect 13486 24652 13492 24654
rect 13556 24652 13562 24716
rect 13997 24714 14063 24717
rect 13997 24712 14842 24714
rect 13997 24656 14002 24712
rect 14058 24656 14842 24712
rect 13997 24654 14842 24656
rect 13997 24651 14063 24654
rect 0 24578 160 24608
rect 749 24578 815 24581
rect 0 24576 815 24578
rect 0 24520 754 24576
rect 810 24520 815 24576
rect 0 24518 815 24520
rect 14782 24578 14842 24654
rect 15840 24578 16000 24608
rect 14782 24518 16000 24578
rect 0 24488 160 24518
rect 749 24515 815 24518
rect 2659 24512 2975 24513
rect 2659 24448 2665 24512
rect 2729 24448 2745 24512
rect 2809 24448 2825 24512
rect 2889 24448 2905 24512
rect 2969 24448 2975 24512
rect 2659 24447 2975 24448
rect 6086 24512 6402 24513
rect 6086 24448 6092 24512
rect 6156 24448 6172 24512
rect 6236 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6402 24512
rect 6086 24447 6402 24448
rect 9513 24512 9829 24513
rect 9513 24448 9519 24512
rect 9583 24448 9599 24512
rect 9663 24448 9679 24512
rect 9743 24448 9759 24512
rect 9823 24448 9829 24512
rect 9513 24447 9829 24448
rect 12940 24512 13256 24513
rect 12940 24448 12946 24512
rect 13010 24448 13026 24512
rect 13090 24448 13106 24512
rect 13170 24448 13186 24512
rect 13250 24448 13256 24512
rect 15840 24488 16000 24518
rect 12940 24447 13256 24448
rect 5901 24306 5967 24309
rect 8661 24306 8727 24309
rect 9489 24306 9555 24309
rect 5901 24304 9555 24306
rect 5901 24248 5906 24304
rect 5962 24248 8666 24304
rect 8722 24248 9494 24304
rect 9550 24248 9555 24304
rect 5901 24246 9555 24248
rect 5901 24243 5967 24246
rect 8661 24243 8727 24246
rect 9489 24243 9555 24246
rect 11973 24306 12039 24309
rect 15840 24306 16000 24336
rect 11973 24304 16000 24306
rect 11973 24248 11978 24304
rect 12034 24248 16000 24304
rect 11973 24246 16000 24248
rect 11973 24243 12039 24246
rect 15840 24216 16000 24246
rect 13905 24170 13971 24173
rect 13905 24168 14474 24170
rect 13905 24112 13910 24168
rect 13966 24112 14474 24168
rect 13905 24110 14474 24112
rect 13905 24107 13971 24110
rect 7189 24034 7255 24037
rect 7414 24034 7420 24036
rect 7189 24032 7420 24034
rect 7189 23976 7194 24032
rect 7250 23976 7420 24032
rect 7189 23974 7420 23976
rect 7189 23971 7255 23974
rect 7414 23972 7420 23974
rect 7484 23972 7490 24036
rect 4372 23968 4688 23969
rect 4372 23904 4378 23968
rect 4442 23904 4458 23968
rect 4522 23904 4538 23968
rect 4602 23904 4618 23968
rect 4682 23904 4688 23968
rect 4372 23903 4688 23904
rect 7799 23968 8115 23969
rect 7799 23904 7805 23968
rect 7869 23904 7885 23968
rect 7949 23904 7965 23968
rect 8029 23904 8045 23968
rect 8109 23904 8115 23968
rect 7799 23903 8115 23904
rect 11226 23968 11542 23969
rect 11226 23904 11232 23968
rect 11296 23904 11312 23968
rect 11376 23904 11392 23968
rect 11456 23904 11472 23968
rect 11536 23904 11542 23968
rect 11226 23903 11542 23904
rect 7097 23898 7163 23901
rect 7414 23898 7420 23900
rect 7097 23896 7420 23898
rect 7097 23840 7102 23896
rect 7158 23840 7420 23896
rect 7097 23838 7420 23840
rect 7097 23835 7163 23838
rect 7414 23836 7420 23838
rect 7484 23836 7490 23900
rect 0 23762 160 23792
rect 749 23762 815 23765
rect 0 23760 815 23762
rect 0 23704 754 23760
rect 810 23704 815 23760
rect 0 23702 815 23704
rect 14414 23762 14474 24110
rect 15101 24034 15167 24037
rect 15840 24034 16000 24064
rect 15101 24032 16000 24034
rect 15101 23976 15106 24032
rect 15162 23976 16000 24032
rect 15101 23974 16000 23976
rect 15101 23971 15167 23974
rect 14653 23968 14969 23969
rect 14653 23904 14659 23968
rect 14723 23904 14739 23968
rect 14803 23904 14819 23968
rect 14883 23904 14899 23968
rect 14963 23904 14969 23968
rect 15840 23944 16000 23974
rect 14653 23903 14969 23904
rect 15840 23762 16000 23792
rect 14414 23702 16000 23762
rect 0 23672 160 23702
rect 749 23699 815 23702
rect 15840 23672 16000 23702
rect 14181 23490 14247 23493
rect 15840 23490 16000 23520
rect 14181 23488 16000 23490
rect 14181 23432 14186 23488
rect 14242 23432 16000 23488
rect 14181 23430 16000 23432
rect 14181 23427 14247 23430
rect 2659 23424 2975 23425
rect 2659 23360 2665 23424
rect 2729 23360 2745 23424
rect 2809 23360 2825 23424
rect 2889 23360 2905 23424
rect 2969 23360 2975 23424
rect 2659 23359 2975 23360
rect 6086 23424 6402 23425
rect 6086 23360 6092 23424
rect 6156 23360 6172 23424
rect 6236 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6402 23424
rect 6086 23359 6402 23360
rect 9513 23424 9829 23425
rect 9513 23360 9519 23424
rect 9583 23360 9599 23424
rect 9663 23360 9679 23424
rect 9743 23360 9759 23424
rect 9823 23360 9829 23424
rect 9513 23359 9829 23360
rect 12940 23424 13256 23425
rect 12940 23360 12946 23424
rect 13010 23360 13026 23424
rect 13090 23360 13106 23424
rect 13170 23360 13186 23424
rect 13250 23360 13256 23424
rect 15840 23400 16000 23430
rect 12940 23359 13256 23360
rect 1669 23218 1735 23221
rect 7230 23218 7236 23220
rect 1669 23216 7236 23218
rect 1669 23160 1674 23216
rect 1730 23160 7236 23216
rect 1669 23158 7236 23160
rect 1669 23155 1735 23158
rect 7230 23156 7236 23158
rect 7300 23156 7306 23220
rect 14365 23218 14431 23221
rect 15840 23218 16000 23248
rect 14365 23216 16000 23218
rect 14365 23160 14370 23216
rect 14426 23160 16000 23216
rect 14365 23158 16000 23160
rect 14365 23155 14431 23158
rect 15840 23128 16000 23158
rect 8845 23084 8911 23085
rect 12617 23084 12683 23085
rect 8845 23082 8892 23084
rect 8804 23080 8892 23082
rect 8956 23082 8962 23084
rect 11646 23082 11652 23084
rect 8804 23024 8850 23080
rect 8804 23022 8892 23024
rect 8845 23020 8892 23022
rect 8956 23022 11652 23082
rect 8956 23020 8962 23022
rect 11646 23020 11652 23022
rect 11716 23020 11722 23084
rect 12566 23020 12572 23084
rect 12636 23082 12683 23084
rect 12636 23080 12728 23082
rect 12678 23024 12728 23080
rect 12636 23022 12728 23024
rect 12636 23020 12683 23022
rect 8845 23019 8911 23020
rect 12617 23019 12683 23020
rect 0 22946 160 22976
rect 749 22946 815 22949
rect 0 22944 815 22946
rect 0 22888 754 22944
rect 810 22888 815 22944
rect 0 22886 815 22888
rect 0 22856 160 22886
rect 749 22883 815 22886
rect 15101 22946 15167 22949
rect 15840 22946 16000 22976
rect 15101 22944 16000 22946
rect 15101 22888 15106 22944
rect 15162 22888 16000 22944
rect 15101 22886 16000 22888
rect 15101 22883 15167 22886
rect 4372 22880 4688 22881
rect 4372 22816 4378 22880
rect 4442 22816 4458 22880
rect 4522 22816 4538 22880
rect 4602 22816 4618 22880
rect 4682 22816 4688 22880
rect 4372 22815 4688 22816
rect 7799 22880 8115 22881
rect 7799 22816 7805 22880
rect 7869 22816 7885 22880
rect 7949 22816 7965 22880
rect 8029 22816 8045 22880
rect 8109 22816 8115 22880
rect 7799 22815 8115 22816
rect 11226 22880 11542 22881
rect 11226 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11392 22880
rect 11456 22816 11472 22880
rect 11536 22816 11542 22880
rect 11226 22815 11542 22816
rect 14653 22880 14969 22881
rect 14653 22816 14659 22880
rect 14723 22816 14739 22880
rect 14803 22816 14819 22880
rect 14883 22816 14899 22880
rect 14963 22816 14969 22880
rect 15840 22856 16000 22886
rect 14653 22815 14969 22816
rect 8385 22674 8451 22677
rect 9254 22674 9260 22676
rect 8385 22672 9260 22674
rect 8385 22616 8390 22672
rect 8446 22616 9260 22672
rect 8385 22614 9260 22616
rect 8385 22611 8451 22614
rect 9254 22612 9260 22614
rect 9324 22612 9330 22676
rect 11145 22674 11211 22677
rect 11830 22674 11836 22676
rect 11145 22672 11836 22674
rect 11145 22616 11150 22672
rect 11206 22616 11836 22672
rect 11145 22614 11836 22616
rect 11145 22611 11211 22614
rect 11830 22612 11836 22614
rect 11900 22612 11906 22676
rect 14273 22674 14339 22677
rect 15840 22674 16000 22704
rect 14273 22672 16000 22674
rect 14273 22616 14278 22672
rect 14334 22616 16000 22672
rect 14273 22614 16000 22616
rect 14273 22611 14339 22614
rect 15840 22584 16000 22614
rect 8886 22476 8892 22540
rect 8956 22538 8962 22540
rect 13537 22538 13603 22541
rect 8956 22536 13603 22538
rect 8956 22480 13542 22536
rect 13598 22480 13603 22536
rect 8956 22478 13603 22480
rect 8956 22476 8962 22478
rect 13537 22475 13603 22478
rect 13721 22402 13787 22405
rect 15840 22402 16000 22432
rect 13721 22400 16000 22402
rect 13721 22344 13726 22400
rect 13782 22344 16000 22400
rect 13721 22342 16000 22344
rect 13721 22339 13787 22342
rect 2659 22336 2975 22337
rect 2659 22272 2665 22336
rect 2729 22272 2745 22336
rect 2809 22272 2825 22336
rect 2889 22272 2905 22336
rect 2969 22272 2975 22336
rect 2659 22271 2975 22272
rect 6086 22336 6402 22337
rect 6086 22272 6092 22336
rect 6156 22272 6172 22336
rect 6236 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6402 22336
rect 6086 22271 6402 22272
rect 9513 22336 9829 22337
rect 9513 22272 9519 22336
rect 9583 22272 9599 22336
rect 9663 22272 9679 22336
rect 9743 22272 9759 22336
rect 9823 22272 9829 22336
rect 9513 22271 9829 22272
rect 12940 22336 13256 22337
rect 12940 22272 12946 22336
rect 13010 22272 13026 22336
rect 13090 22272 13106 22336
rect 13170 22272 13186 22336
rect 13250 22272 13256 22336
rect 15840 22312 16000 22342
rect 12940 22271 13256 22272
rect 0 22130 160 22160
rect 749 22130 815 22133
rect 0 22128 815 22130
rect 0 22072 754 22128
rect 810 22072 815 22128
rect 0 22070 815 22072
rect 0 22040 160 22070
rect 749 22067 815 22070
rect 12157 22130 12223 22133
rect 12750 22130 12756 22132
rect 12157 22128 12756 22130
rect 12157 22072 12162 22128
rect 12218 22072 12756 22128
rect 12157 22070 12756 22072
rect 12157 22067 12223 22070
rect 12750 22068 12756 22070
rect 12820 22068 12826 22132
rect 13813 22130 13879 22133
rect 15840 22130 16000 22160
rect 13813 22128 16000 22130
rect 13813 22072 13818 22128
rect 13874 22072 16000 22128
rect 13813 22070 16000 22072
rect 13813 22067 13879 22070
rect 15840 22040 16000 22070
rect 7557 21996 7623 21997
rect 7557 21994 7604 21996
rect 7512 21992 7604 21994
rect 7512 21936 7562 21992
rect 7512 21934 7604 21936
rect 7557 21932 7604 21934
rect 7668 21932 7674 21996
rect 9857 21994 9923 21997
rect 14365 21994 14431 21997
rect 9857 21992 14431 21994
rect 9857 21936 9862 21992
rect 9918 21936 14370 21992
rect 14426 21936 14431 21992
rect 9857 21934 14431 21936
rect 7557 21931 7623 21932
rect 9857 21931 9923 21934
rect 14365 21931 14431 21934
rect 15193 21858 15259 21861
rect 15840 21858 16000 21888
rect 15193 21856 16000 21858
rect 15193 21800 15198 21856
rect 15254 21800 16000 21856
rect 15193 21798 16000 21800
rect 15193 21795 15259 21798
rect 4372 21792 4688 21793
rect 4372 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4688 21792
rect 4372 21727 4688 21728
rect 7799 21792 8115 21793
rect 7799 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8115 21792
rect 7799 21727 8115 21728
rect 11226 21792 11542 21793
rect 11226 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11542 21792
rect 11226 21727 11542 21728
rect 14653 21792 14969 21793
rect 14653 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14969 21792
rect 15840 21768 16000 21798
rect 14653 21727 14969 21728
rect 9765 21722 9831 21725
rect 9990 21722 9996 21724
rect 9765 21720 9996 21722
rect 9765 21664 9770 21720
rect 9826 21664 9996 21720
rect 9765 21662 9996 21664
rect 9765 21659 9831 21662
rect 9990 21660 9996 21662
rect 10060 21660 10066 21724
rect 6269 21586 6335 21589
rect 12801 21586 12867 21589
rect 13629 21586 13695 21589
rect 6269 21584 13695 21586
rect 6269 21528 6274 21584
rect 6330 21528 12806 21584
rect 12862 21528 13634 21584
rect 13690 21528 13695 21584
rect 6269 21526 13695 21528
rect 6269 21523 6335 21526
rect 12801 21523 12867 21526
rect 13629 21523 13695 21526
rect 14089 21586 14155 21589
rect 15840 21586 16000 21616
rect 14089 21584 16000 21586
rect 14089 21528 14094 21584
rect 14150 21528 16000 21584
rect 14089 21526 16000 21528
rect 14089 21523 14155 21526
rect 15840 21496 16000 21526
rect 11789 21450 11855 21453
rect 11789 21448 14290 21450
rect 11789 21392 11794 21448
rect 11850 21392 14290 21448
rect 11789 21390 14290 21392
rect 11789 21387 11855 21390
rect 0 21314 160 21344
rect 749 21314 815 21317
rect 0 21312 815 21314
rect 0 21256 754 21312
rect 810 21256 815 21312
rect 0 21254 815 21256
rect 14230 21314 14290 21390
rect 15840 21314 16000 21344
rect 14230 21254 16000 21314
rect 0 21224 160 21254
rect 749 21251 815 21254
rect 2659 21248 2975 21249
rect 2659 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2975 21248
rect 2659 21183 2975 21184
rect 6086 21248 6402 21249
rect 6086 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6402 21248
rect 6086 21183 6402 21184
rect 9513 21248 9829 21249
rect 9513 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9829 21248
rect 9513 21183 9829 21184
rect 12940 21248 13256 21249
rect 12940 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13256 21248
rect 15840 21224 16000 21254
rect 12940 21183 13256 21184
rect 12249 21180 12315 21181
rect 12198 21116 12204 21180
rect 12268 21178 12315 21180
rect 12268 21176 12360 21178
rect 12310 21120 12360 21176
rect 12268 21118 12360 21120
rect 12268 21116 12315 21118
rect 12249 21115 12315 21116
rect 12157 21042 12223 21045
rect 13905 21042 13971 21045
rect 12157 21040 13971 21042
rect 12157 20984 12162 21040
rect 12218 20984 13910 21040
rect 13966 20984 13971 21040
rect 12157 20982 13971 20984
rect 12157 20979 12223 20982
rect 13905 20979 13971 20982
rect 14273 21042 14339 21045
rect 15840 21042 16000 21072
rect 14273 21040 16000 21042
rect 14273 20984 14278 21040
rect 14334 20984 16000 21040
rect 14273 20982 16000 20984
rect 14273 20979 14339 20982
rect 15840 20952 16000 20982
rect 7005 20906 7071 20909
rect 8937 20906 9003 20909
rect 7005 20904 9003 20906
rect 7005 20848 7010 20904
rect 7066 20848 8942 20904
rect 8998 20848 9003 20904
rect 7005 20846 9003 20848
rect 7005 20843 7071 20846
rect 8937 20843 9003 20846
rect 11973 20906 12039 20909
rect 11973 20904 15210 20906
rect 11973 20848 11978 20904
rect 12034 20848 15210 20904
rect 11973 20846 15210 20848
rect 11973 20843 12039 20846
rect 15150 20770 15210 20846
rect 15840 20770 16000 20800
rect 15150 20710 16000 20770
rect 4372 20704 4688 20705
rect 4372 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4688 20704
rect 4372 20639 4688 20640
rect 7799 20704 8115 20705
rect 7799 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8115 20704
rect 7799 20639 8115 20640
rect 11226 20704 11542 20705
rect 11226 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11542 20704
rect 11226 20639 11542 20640
rect 14653 20704 14969 20705
rect 14653 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14969 20704
rect 15840 20680 16000 20710
rect 14653 20639 14969 20640
rect 1393 20634 1459 20637
rect 752 20632 1459 20634
rect 752 20576 1398 20632
rect 1454 20576 1459 20632
rect 752 20574 1459 20576
rect 0 20498 160 20528
rect 752 20498 812 20574
rect 1393 20571 1459 20574
rect 0 20438 812 20498
rect 12525 20498 12591 20501
rect 15840 20498 16000 20528
rect 12525 20496 16000 20498
rect 12525 20440 12530 20496
rect 12586 20440 16000 20496
rect 12525 20438 16000 20440
rect 0 20408 160 20438
rect 12525 20435 12591 20438
rect 15840 20408 16000 20438
rect 1945 20362 2011 20365
rect 11053 20362 11119 20365
rect 12341 20362 12407 20365
rect 1945 20360 12407 20362
rect 1945 20304 1950 20360
rect 2006 20304 11058 20360
rect 11114 20304 12346 20360
rect 12402 20304 12407 20360
rect 1945 20302 12407 20304
rect 1945 20299 2011 20302
rect 11053 20299 11119 20302
rect 12341 20299 12407 20302
rect 14365 20226 14431 20229
rect 15840 20226 16000 20256
rect 14365 20224 16000 20226
rect 14365 20168 14370 20224
rect 14426 20168 16000 20224
rect 14365 20166 16000 20168
rect 14365 20163 14431 20166
rect 2659 20160 2975 20161
rect 2659 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2975 20160
rect 2659 20095 2975 20096
rect 6086 20160 6402 20161
rect 6086 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6402 20160
rect 6086 20095 6402 20096
rect 9513 20160 9829 20161
rect 9513 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9829 20160
rect 9513 20095 9829 20096
rect 12940 20160 13256 20161
rect 12940 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13256 20160
rect 15840 20136 16000 20166
rect 12940 20095 13256 20096
rect 9949 20090 10015 20093
rect 9949 20088 10058 20090
rect 9949 20032 9954 20088
rect 10010 20032 10058 20088
rect 9949 20027 10058 20032
rect 10133 20088 10199 20093
rect 10133 20032 10138 20088
rect 10194 20032 10199 20088
rect 10133 20027 10199 20032
rect 9998 19954 10058 20027
rect 9860 19894 10058 19954
rect 0 19682 160 19712
rect 9860 19685 9920 19894
rect 10136 19685 10196 20027
rect 13077 19954 13143 19957
rect 13670 19954 13676 19956
rect 13077 19952 13676 19954
rect 13077 19896 13082 19952
rect 13138 19896 13676 19952
rect 13077 19894 13676 19896
rect 13077 19891 13143 19894
rect 13670 19892 13676 19894
rect 13740 19892 13746 19956
rect 13905 19954 13971 19957
rect 15840 19954 16000 19984
rect 13905 19952 16000 19954
rect 13905 19896 13910 19952
rect 13966 19896 16000 19952
rect 13905 19894 16000 19896
rect 13905 19891 13971 19894
rect 15840 19864 16000 19894
rect 749 19682 815 19685
rect 0 19680 815 19682
rect 0 19624 754 19680
rect 810 19624 815 19680
rect 0 19622 815 19624
rect 0 19592 160 19622
rect 749 19619 815 19622
rect 9857 19680 9923 19685
rect 9857 19624 9862 19680
rect 9918 19624 9923 19680
rect 9857 19619 9923 19624
rect 10133 19680 10199 19685
rect 10133 19624 10138 19680
rect 10194 19624 10199 19680
rect 10133 19619 10199 19624
rect 15469 19682 15535 19685
rect 15840 19682 16000 19712
rect 15469 19680 16000 19682
rect 15469 19624 15474 19680
rect 15530 19624 16000 19680
rect 15469 19622 16000 19624
rect 15469 19619 15535 19622
rect 4372 19616 4688 19617
rect 4372 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4688 19616
rect 4372 19551 4688 19552
rect 7799 19616 8115 19617
rect 7799 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8115 19616
rect 7799 19551 8115 19552
rect 11226 19616 11542 19617
rect 11226 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11542 19616
rect 11226 19551 11542 19552
rect 14653 19616 14969 19617
rect 14653 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14969 19616
rect 15840 19592 16000 19622
rect 14653 19551 14969 19552
rect 9029 19548 9095 19549
rect 10041 19548 10107 19549
rect 9029 19544 9076 19548
rect 9140 19546 9146 19548
rect 9990 19546 9996 19548
rect 9029 19488 9034 19544
rect 9029 19484 9076 19488
rect 9140 19486 9186 19546
rect 9950 19486 9996 19546
rect 10060 19544 10107 19548
rect 10102 19488 10107 19544
rect 9140 19484 9146 19486
rect 9990 19484 9996 19486
rect 10060 19484 10107 19488
rect 9029 19483 9095 19484
rect 10041 19483 10107 19484
rect 5533 19410 5599 19413
rect 10961 19410 11027 19413
rect 5533 19408 11027 19410
rect 5533 19352 5538 19408
rect 5594 19352 10966 19408
rect 11022 19352 11027 19408
rect 5533 19350 11027 19352
rect 5533 19347 5599 19350
rect 10961 19347 11027 19350
rect 13813 19410 13879 19413
rect 15840 19410 16000 19440
rect 13813 19408 16000 19410
rect 13813 19352 13818 19408
rect 13874 19352 16000 19408
rect 13813 19350 16000 19352
rect 13813 19347 13879 19350
rect 15840 19320 16000 19350
rect 1485 19272 1551 19277
rect 1485 19216 1490 19272
rect 1546 19216 1551 19272
rect 1485 19211 1551 19216
rect 1669 19274 1735 19277
rect 1669 19272 11898 19274
rect 1669 19216 1674 19272
rect 1730 19216 11898 19272
rect 1669 19214 11898 19216
rect 1669 19211 1735 19214
rect 0 18866 160 18896
rect 1488 18866 1548 19211
rect 2659 19072 2975 19073
rect 2659 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2975 19072
rect 2659 19007 2975 19008
rect 6086 19072 6402 19073
rect 6086 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6402 19072
rect 6086 19007 6402 19008
rect 9513 19072 9829 19073
rect 9513 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9829 19072
rect 9513 19007 9829 19008
rect 7833 19002 7899 19005
rect 11838 19004 11898 19214
rect 14273 19138 14339 19141
rect 15840 19138 16000 19168
rect 14273 19136 16000 19138
rect 14273 19080 14278 19136
rect 14334 19080 16000 19136
rect 14273 19078 16000 19080
rect 14273 19075 14339 19078
rect 12940 19072 13256 19073
rect 12940 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13256 19072
rect 15840 19048 16000 19078
rect 12940 19007 13256 19008
rect 7238 19000 7899 19002
rect 7238 18944 7838 19000
rect 7894 18944 7899 19000
rect 7238 18942 7899 18944
rect 0 18806 1548 18866
rect 3509 18866 3575 18869
rect 7238 18866 7298 18942
rect 7833 18939 7899 18942
rect 11830 18940 11836 19004
rect 11900 19002 11906 19004
rect 11900 18942 12772 19002
rect 11900 18940 11906 18942
rect 3509 18864 7298 18866
rect 3509 18808 3514 18864
rect 3570 18808 7298 18864
rect 3509 18806 7298 18808
rect 7373 18868 7439 18869
rect 7373 18864 7420 18868
rect 7484 18866 7490 18868
rect 9581 18866 9647 18869
rect 12566 18866 12572 18868
rect 7373 18808 7378 18864
rect 0 18776 160 18806
rect 3509 18803 3575 18806
rect 7373 18804 7420 18808
rect 7484 18806 7530 18866
rect 9581 18864 12572 18866
rect 9581 18808 9586 18864
rect 9642 18808 12572 18864
rect 9581 18806 12572 18808
rect 7484 18804 7490 18806
rect 7373 18803 7439 18804
rect 9581 18803 9647 18806
rect 12566 18804 12572 18806
rect 12636 18804 12642 18868
rect 12712 18866 12772 18942
rect 12985 18866 13051 18869
rect 12712 18864 13051 18866
rect 12712 18808 12990 18864
rect 13046 18808 13051 18864
rect 12712 18806 13051 18808
rect 12985 18803 13051 18806
rect 14089 18866 14155 18869
rect 15840 18866 16000 18896
rect 14089 18864 16000 18866
rect 14089 18808 14094 18864
rect 14150 18808 16000 18864
rect 14089 18806 16000 18808
rect 14089 18803 14155 18806
rect 15840 18776 16000 18806
rect 7414 18668 7420 18732
rect 7484 18730 7490 18732
rect 7649 18730 7715 18733
rect 7484 18728 7715 18730
rect 7484 18672 7654 18728
rect 7710 18672 7715 18728
rect 7484 18670 7715 18672
rect 7484 18668 7490 18670
rect 7649 18667 7715 18670
rect 9673 18730 9739 18733
rect 10726 18730 10732 18732
rect 9673 18728 10732 18730
rect 9673 18672 9678 18728
rect 9734 18672 10732 18728
rect 9673 18670 10732 18672
rect 9673 18667 9739 18670
rect 10726 18668 10732 18670
rect 10796 18668 10802 18732
rect 11789 18730 11855 18733
rect 11789 18728 15578 18730
rect 11789 18672 11794 18728
rect 11850 18672 15578 18728
rect 11789 18670 15578 18672
rect 11789 18667 11855 18670
rect 11789 18594 11855 18597
rect 13905 18594 13971 18597
rect 11789 18592 13971 18594
rect 11789 18536 11794 18592
rect 11850 18536 13910 18592
rect 13966 18536 13971 18592
rect 11789 18534 13971 18536
rect 15518 18594 15578 18670
rect 15840 18594 16000 18624
rect 15518 18534 16000 18594
rect 11789 18531 11855 18534
rect 13905 18531 13971 18534
rect 4372 18528 4688 18529
rect 4372 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4688 18528
rect 4372 18463 4688 18464
rect 7799 18528 8115 18529
rect 7799 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8115 18528
rect 7799 18463 8115 18464
rect 11226 18528 11542 18529
rect 11226 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11542 18528
rect 11226 18463 11542 18464
rect 14653 18528 14969 18529
rect 14653 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14969 18528
rect 15840 18504 16000 18534
rect 14653 18463 14969 18464
rect 13905 18322 13971 18325
rect 15840 18322 16000 18352
rect 13905 18320 16000 18322
rect 13905 18264 13910 18320
rect 13966 18264 16000 18320
rect 13905 18262 16000 18264
rect 13905 18259 13971 18262
rect 15840 18232 16000 18262
rect 11421 18186 11487 18189
rect 11421 18184 14290 18186
rect 11421 18128 11426 18184
rect 11482 18128 14290 18184
rect 11421 18126 14290 18128
rect 11421 18123 11487 18126
rect 0 18050 160 18080
rect 749 18050 815 18053
rect 0 18048 815 18050
rect 0 17992 754 18048
rect 810 17992 815 18048
rect 0 17990 815 17992
rect 0 17960 160 17990
rect 749 17987 815 17990
rect 10133 18050 10199 18053
rect 12433 18050 12499 18053
rect 10133 18048 12499 18050
rect 10133 17992 10138 18048
rect 10194 17992 12438 18048
rect 12494 17992 12499 18048
rect 10133 17990 12499 17992
rect 14230 18050 14290 18126
rect 15840 18050 16000 18080
rect 14230 17990 16000 18050
rect 10133 17987 10199 17990
rect 12433 17987 12499 17990
rect 2659 17984 2975 17985
rect 2659 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2975 17984
rect 2659 17919 2975 17920
rect 6086 17984 6402 17985
rect 6086 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6402 17984
rect 6086 17919 6402 17920
rect 9513 17984 9829 17985
rect 9513 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9829 17984
rect 9513 17919 9829 17920
rect 12940 17984 13256 17985
rect 12940 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13256 17984
rect 15840 17960 16000 17990
rect 12940 17919 13256 17920
rect 10409 17914 10475 17917
rect 11789 17914 11855 17917
rect 13813 17916 13879 17917
rect 13813 17914 13860 17916
rect 10409 17912 11855 17914
rect 10409 17856 10414 17912
rect 10470 17856 11794 17912
rect 11850 17856 11855 17912
rect 10409 17854 11855 17856
rect 13768 17912 13860 17914
rect 13768 17856 13818 17912
rect 13768 17854 13860 17856
rect 10409 17851 10475 17854
rect 11789 17851 11855 17854
rect 13813 17852 13860 17854
rect 13924 17852 13930 17916
rect 14549 17914 14615 17917
rect 15193 17914 15259 17917
rect 14549 17912 15259 17914
rect 14549 17856 14554 17912
rect 14610 17856 15198 17912
rect 15254 17856 15259 17912
rect 14549 17854 15259 17856
rect 13813 17851 13879 17852
rect 14549 17851 14615 17854
rect 15193 17851 15259 17854
rect 5441 17778 5507 17781
rect 9673 17778 9739 17781
rect 10542 17778 10548 17780
rect 5441 17776 6746 17778
rect 5441 17720 5446 17776
rect 5502 17720 6746 17776
rect 5441 17718 6746 17720
rect 5441 17715 5507 17718
rect 6453 17644 6519 17645
rect 6453 17640 6500 17644
rect 6564 17642 6570 17644
rect 6686 17642 6746 17718
rect 9673 17776 10548 17778
rect 9673 17720 9678 17776
rect 9734 17720 10548 17776
rect 9673 17718 10548 17720
rect 9673 17715 9739 17718
rect 10542 17716 10548 17718
rect 10612 17716 10618 17780
rect 11145 17778 11211 17781
rect 15840 17778 16000 17808
rect 11145 17776 16000 17778
rect 11145 17720 11150 17776
rect 11206 17720 16000 17776
rect 11145 17718 16000 17720
rect 11145 17715 11211 17718
rect 15840 17688 16000 17718
rect 11830 17642 11836 17644
rect 6453 17584 6458 17640
rect 6453 17580 6500 17584
rect 6564 17582 6610 17642
rect 6686 17582 11836 17642
rect 6564 17580 6570 17582
rect 11830 17580 11836 17582
rect 11900 17580 11906 17644
rect 6453 17579 6519 17580
rect 11789 17506 11855 17509
rect 13721 17506 13787 17509
rect 11789 17504 13787 17506
rect 11789 17448 11794 17504
rect 11850 17448 13726 17504
rect 13782 17448 13787 17504
rect 11789 17446 13787 17448
rect 11789 17443 11855 17446
rect 13721 17443 13787 17446
rect 14181 17508 14247 17509
rect 14181 17504 14228 17508
rect 14292 17506 14298 17508
rect 15193 17506 15259 17509
rect 15840 17506 16000 17536
rect 14181 17448 14186 17504
rect 14181 17444 14228 17448
rect 14292 17446 14338 17506
rect 15193 17504 16000 17506
rect 15193 17448 15198 17504
rect 15254 17448 16000 17504
rect 15193 17446 16000 17448
rect 14292 17444 14298 17446
rect 14181 17443 14247 17444
rect 15193 17443 15259 17446
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 15840 17416 16000 17446
rect 14653 17375 14969 17376
rect 12525 17370 12591 17373
rect 13486 17370 13492 17372
rect 12525 17368 13492 17370
rect 12525 17312 12530 17368
rect 12586 17312 13492 17368
rect 12525 17310 13492 17312
rect 12525 17307 12591 17310
rect 13486 17308 13492 17310
rect 13556 17308 13562 17372
rect 0 17234 160 17264
rect 749 17234 815 17237
rect 0 17232 815 17234
rect 0 17176 754 17232
rect 810 17176 815 17232
rect 0 17174 815 17176
rect 0 17144 160 17174
rect 749 17171 815 17174
rect 11697 17234 11763 17237
rect 15840 17234 16000 17264
rect 11697 17232 16000 17234
rect 11697 17176 11702 17232
rect 11758 17176 16000 17232
rect 11697 17174 16000 17176
rect 11697 17171 11763 17174
rect 15840 17144 16000 17174
rect 5165 17098 5231 17101
rect 9673 17098 9739 17101
rect 5165 17096 9739 17098
rect 5165 17040 5170 17096
rect 5226 17040 9678 17096
rect 9734 17040 9739 17096
rect 5165 17038 9739 17040
rect 5165 17035 5231 17038
rect 9673 17035 9739 17038
rect 11421 17098 11487 17101
rect 11646 17098 11652 17100
rect 11421 17096 11652 17098
rect 11421 17040 11426 17096
rect 11482 17040 11652 17096
rect 11421 17038 11652 17040
rect 11421 17035 11487 17038
rect 11646 17036 11652 17038
rect 11716 17036 11722 17100
rect 11789 17098 11855 17101
rect 14549 17098 14615 17101
rect 11789 17096 14615 17098
rect 11789 17040 11794 17096
rect 11850 17040 14554 17096
rect 14610 17040 14615 17096
rect 11789 17038 14615 17040
rect 11654 16962 11714 17036
rect 11789 17035 11855 17038
rect 14549 17035 14615 17038
rect 12065 16962 12131 16965
rect 11654 16960 12131 16962
rect 11654 16904 12070 16960
rect 12126 16904 12131 16960
rect 11654 16902 12131 16904
rect 12065 16899 12131 16902
rect 14549 16962 14615 16965
rect 15840 16962 16000 16992
rect 14549 16960 16000 16962
rect 14549 16904 14554 16960
rect 14610 16904 16000 16960
rect 14549 16902 16000 16904
rect 14549 16899 14615 16902
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 15840 16872 16000 16902
rect 12940 16831 13256 16832
rect 10133 16826 10199 16829
rect 12198 16826 12204 16828
rect 10133 16824 12204 16826
rect 10133 16768 10138 16824
rect 10194 16768 12204 16824
rect 10133 16766 12204 16768
rect 10133 16763 10199 16766
rect 12198 16764 12204 16766
rect 12268 16826 12274 16828
rect 12525 16826 12591 16829
rect 12268 16824 12591 16826
rect 12268 16768 12530 16824
rect 12586 16768 12591 16824
rect 12268 16766 12591 16768
rect 12268 16764 12274 16766
rect 12525 16763 12591 16766
rect 12893 16690 12959 16693
rect 14038 16690 14044 16692
rect 12893 16688 14044 16690
rect 12893 16632 12898 16688
rect 12954 16632 14044 16688
rect 12893 16630 14044 16632
rect 12893 16627 12959 16630
rect 14038 16628 14044 16630
rect 14108 16628 14114 16692
rect 14273 16690 14339 16693
rect 15840 16690 16000 16720
rect 14273 16688 16000 16690
rect 14273 16632 14278 16688
rect 14334 16632 16000 16688
rect 14273 16630 16000 16632
rect 14273 16627 14339 16630
rect 15840 16600 16000 16630
rect 1485 16554 1551 16557
rect 798 16552 1551 16554
rect 798 16496 1490 16552
rect 1546 16496 1551 16552
rect 798 16494 1551 16496
rect 0 16418 160 16448
rect 798 16418 858 16494
rect 1485 16491 1551 16494
rect 7557 16556 7623 16557
rect 9213 16556 9279 16557
rect 7557 16552 7604 16556
rect 7668 16554 7674 16556
rect 9213 16554 9260 16556
rect 7557 16496 7562 16552
rect 7557 16492 7604 16496
rect 7668 16494 7714 16554
rect 9168 16552 9260 16554
rect 9168 16496 9218 16552
rect 9168 16494 9260 16496
rect 7668 16492 7674 16494
rect 9213 16492 9260 16494
rect 9324 16492 9330 16556
rect 13724 16494 15210 16554
rect 7557 16491 7623 16492
rect 9213 16491 9279 16492
rect 13724 16421 13784 16494
rect 0 16358 858 16418
rect 9949 16418 10015 16421
rect 10542 16418 10548 16420
rect 9949 16416 10548 16418
rect 9949 16360 9954 16416
rect 10010 16360 10548 16416
rect 9949 16358 10548 16360
rect 0 16328 160 16358
rect 9949 16355 10015 16358
rect 10542 16356 10548 16358
rect 10612 16356 10618 16420
rect 13721 16416 13787 16421
rect 13721 16360 13726 16416
rect 13782 16360 13787 16416
rect 13721 16355 13787 16360
rect 14181 16416 14247 16421
rect 14181 16360 14186 16416
rect 14242 16360 14247 16416
rect 14181 16355 14247 16360
rect 15150 16418 15210 16494
rect 15840 16418 16000 16448
rect 15150 16358 16000 16418
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14184 16282 14244 16355
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 15840 16328 16000 16358
rect 14653 16287 14969 16288
rect 11884 16222 14244 16282
rect 8937 16146 9003 16149
rect 9305 16146 9371 16149
rect 11884 16146 11944 16222
rect 8937 16144 9138 16146
rect 8937 16088 8942 16144
rect 8998 16088 9138 16144
rect 8937 16086 9138 16088
rect 8937 16083 9003 16086
rect 9078 16010 9138 16086
rect 9305 16144 11944 16146
rect 9305 16088 9310 16144
rect 9366 16088 11944 16144
rect 9305 16086 11944 16088
rect 14181 16146 14247 16149
rect 15840 16146 16000 16176
rect 14181 16144 16000 16146
rect 14181 16088 14186 16144
rect 14242 16088 16000 16144
rect 14181 16086 16000 16088
rect 9305 16083 9371 16086
rect 14181 16083 14247 16086
rect 15840 16056 16000 16086
rect 13445 16010 13511 16013
rect 9078 16008 13511 16010
rect 9078 15952 13450 16008
rect 13506 15952 13511 16008
rect 9078 15950 13511 15952
rect 13445 15947 13511 15950
rect 15653 15874 15719 15877
rect 15840 15874 16000 15904
rect 15653 15872 16000 15874
rect 15653 15816 15658 15872
rect 15714 15816 16000 15872
rect 15653 15814 16000 15816
rect 15653 15811 15719 15814
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 15840 15784 16000 15814
rect 12940 15743 13256 15744
rect 0 15602 160 15632
rect 749 15602 815 15605
rect 0 15600 815 15602
rect 0 15544 754 15600
rect 810 15544 815 15600
rect 0 15542 815 15544
rect 0 15512 160 15542
rect 749 15539 815 15542
rect 13261 15602 13327 15605
rect 15840 15602 16000 15632
rect 13261 15600 16000 15602
rect 13261 15544 13266 15600
rect 13322 15544 16000 15600
rect 13261 15542 16000 15544
rect 13261 15539 13327 15542
rect 15840 15512 16000 15542
rect 14089 15466 14155 15469
rect 14089 15464 15210 15466
rect 14089 15408 14094 15464
rect 14150 15408 15210 15464
rect 14089 15406 15210 15408
rect 14089 15403 14155 15406
rect 12750 15268 12756 15332
rect 12820 15330 12826 15332
rect 14089 15330 14155 15333
rect 12820 15328 14155 15330
rect 12820 15272 14094 15328
rect 14150 15272 14155 15328
rect 12820 15270 14155 15272
rect 15150 15330 15210 15406
rect 15840 15330 16000 15360
rect 15150 15270 16000 15330
rect 12820 15268 12826 15270
rect 14089 15267 14155 15270
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 15840 15240 16000 15270
rect 14653 15199 14969 15200
rect 8201 15194 8267 15197
rect 8886 15194 8892 15196
rect 8201 15192 8892 15194
rect 8201 15136 8206 15192
rect 8262 15136 8892 15192
rect 8201 15134 8892 15136
rect 8201 15131 8267 15134
rect 8886 15132 8892 15134
rect 8956 15132 8962 15196
rect 12750 15132 12756 15196
rect 12820 15194 12826 15196
rect 13077 15194 13143 15197
rect 12820 15192 13143 15194
rect 12820 15136 13082 15192
rect 13138 15136 13143 15192
rect 12820 15134 13143 15136
rect 12820 15132 12826 15134
rect 13077 15131 13143 15134
rect 11973 15058 12039 15061
rect 15840 15058 16000 15088
rect 11973 15056 16000 15058
rect 11973 15000 11978 15056
rect 12034 15000 16000 15056
rect 11973 14998 16000 15000
rect 11973 14995 12039 14998
rect 15840 14968 16000 14998
rect 12985 14922 13051 14925
rect 13670 14922 13676 14924
rect 12985 14920 13676 14922
rect 12985 14864 12990 14920
rect 13046 14864 13676 14920
rect 12985 14862 13676 14864
rect 12985 14859 13051 14862
rect 13670 14860 13676 14862
rect 13740 14860 13746 14924
rect 0 14786 160 14816
rect 841 14786 907 14789
rect 0 14784 907 14786
rect 0 14728 846 14784
rect 902 14728 907 14784
rect 0 14726 907 14728
rect 0 14696 160 14726
rect 841 14723 907 14726
rect 11973 14786 12039 14789
rect 12709 14786 12775 14789
rect 11973 14784 12775 14786
rect 11973 14728 11978 14784
rect 12034 14728 12714 14784
rect 12770 14728 12775 14784
rect 11973 14726 12775 14728
rect 11973 14723 12039 14726
rect 12709 14723 12775 14726
rect 14273 14786 14339 14789
rect 15840 14786 16000 14816
rect 14273 14784 16000 14786
rect 14273 14728 14278 14784
rect 14334 14728 16000 14784
rect 14273 14726 16000 14728
rect 14273 14723 14339 14726
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 15840 14696 16000 14726
rect 12940 14655 13256 14656
rect 11053 14514 11119 14517
rect 11973 14514 12039 14517
rect 11053 14512 12039 14514
rect 11053 14456 11058 14512
rect 11114 14456 11978 14512
rect 12034 14456 12039 14512
rect 11053 14454 12039 14456
rect 11053 14451 11119 14454
rect 11973 14451 12039 14454
rect 15469 14514 15535 14517
rect 15840 14514 16000 14544
rect 15469 14512 16000 14514
rect 15469 14456 15474 14512
rect 15530 14456 16000 14512
rect 15469 14454 16000 14456
rect 15469 14451 15535 14454
rect 15840 14424 16000 14454
rect 7097 14378 7163 14381
rect 7054 14376 7163 14378
rect 7054 14320 7102 14376
rect 7158 14320 7163 14376
rect 7054 14315 7163 14320
rect 10726 14316 10732 14380
rect 10796 14378 10802 14380
rect 10796 14318 11852 14378
rect 10796 14316 10802 14318
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 0 13970 160 14000
rect 841 13970 907 13973
rect 0 13968 907 13970
rect 0 13912 846 13968
rect 902 13912 907 13968
rect 0 13910 907 13912
rect 0 13880 160 13910
rect 841 13907 907 13910
rect 7054 13701 7114 14315
rect 11792 14245 11852 14318
rect 11789 14240 11855 14245
rect 15840 14242 16000 14272
rect 11789 14184 11794 14240
rect 11850 14184 11855 14240
rect 11789 14179 11855 14184
rect 15702 14182 16000 14242
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 14653 14111 14969 14112
rect 15469 14106 15535 14109
rect 15702 14106 15762 14182
rect 15840 14152 16000 14182
rect 15469 14104 15762 14106
rect 15469 14048 15474 14104
rect 15530 14048 15762 14104
rect 15469 14046 15762 14048
rect 15469 14043 15535 14046
rect 9029 13970 9095 13973
rect 9949 13970 10015 13973
rect 12525 13970 12591 13973
rect 9029 13968 12591 13970
rect 9029 13912 9034 13968
rect 9090 13912 9954 13968
rect 10010 13912 12530 13968
rect 12586 13912 12591 13968
rect 9029 13910 12591 13912
rect 9029 13907 9095 13910
rect 9949 13907 10015 13910
rect 12525 13907 12591 13910
rect 13721 13970 13787 13973
rect 15840 13970 16000 14000
rect 13721 13968 16000 13970
rect 13721 13912 13726 13968
rect 13782 13912 16000 13968
rect 13721 13910 16000 13912
rect 13721 13907 13787 13910
rect 15840 13880 16000 13910
rect 10542 13772 10548 13836
rect 10612 13834 10618 13836
rect 11697 13834 11763 13837
rect 14181 13836 14247 13837
rect 14181 13834 14228 13836
rect 10612 13832 11763 13834
rect 10612 13776 11702 13832
rect 11758 13776 11763 13832
rect 10612 13774 11763 13776
rect 14136 13832 14228 13834
rect 14136 13776 14186 13832
rect 14136 13774 14228 13776
rect 10612 13772 10618 13774
rect 11697 13771 11763 13774
rect 14181 13772 14228 13774
rect 14292 13772 14298 13836
rect 14181 13771 14247 13772
rect 7054 13696 7163 13701
rect 7054 13640 7102 13696
rect 7158 13640 7163 13696
rect 7054 13638 7163 13640
rect 7097 13635 7163 13638
rect 14641 13698 14707 13701
rect 15840 13698 16000 13728
rect 14641 13696 16000 13698
rect 14641 13640 14646 13696
rect 14702 13640 16000 13696
rect 14641 13638 16000 13640
rect 14641 13635 14707 13638
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 15840 13608 16000 13638
rect 12940 13567 13256 13568
rect 14181 13426 14247 13429
rect 15840 13426 16000 13456
rect 14181 13424 16000 13426
rect 14181 13368 14186 13424
rect 14242 13368 16000 13424
rect 14181 13366 16000 13368
rect 14181 13363 14247 13366
rect 15840 13336 16000 13366
rect 12249 13290 12315 13293
rect 12617 13290 12683 13293
rect 12249 13288 12683 13290
rect 12249 13232 12254 13288
rect 12310 13232 12622 13288
rect 12678 13232 12683 13288
rect 12249 13230 12683 13232
rect 12249 13227 12315 13230
rect 12617 13227 12683 13230
rect 0 13154 160 13184
rect 841 13154 907 13157
rect 0 13152 907 13154
rect 0 13096 846 13152
rect 902 13096 907 13152
rect 0 13094 907 13096
rect 0 13064 160 13094
rect 841 13091 907 13094
rect 15193 13154 15259 13157
rect 15840 13154 16000 13184
rect 15193 13152 16000 13154
rect 15193 13096 15198 13152
rect 15254 13096 16000 13152
rect 15193 13094 16000 13096
rect 15193 13091 15259 13094
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 15840 13064 16000 13094
rect 14653 13023 14969 13024
rect 7414 12820 7420 12884
rect 7484 12882 7490 12884
rect 8109 12882 8175 12885
rect 7484 12880 8175 12882
rect 7484 12824 8114 12880
rect 8170 12824 8175 12880
rect 7484 12822 8175 12824
rect 7484 12820 7490 12822
rect 8109 12819 8175 12822
rect 12249 12882 12315 12885
rect 13905 12882 13971 12885
rect 12249 12880 13971 12882
rect 12249 12824 12254 12880
rect 12310 12824 13910 12880
rect 13966 12824 13971 12880
rect 12249 12822 13971 12824
rect 12249 12819 12315 12822
rect 13905 12819 13971 12822
rect 14273 12882 14339 12885
rect 15840 12882 16000 12912
rect 14273 12880 16000 12882
rect 14273 12824 14278 12880
rect 14334 12824 16000 12880
rect 14273 12822 16000 12824
rect 14273 12819 14339 12822
rect 15840 12792 16000 12822
rect 3918 12684 3924 12748
rect 3988 12746 3994 12748
rect 14457 12746 14523 12749
rect 3988 12744 14523 12746
rect 3988 12688 14462 12744
rect 14518 12688 14523 12744
rect 3988 12686 14523 12688
rect 3988 12684 3994 12686
rect 14457 12683 14523 12686
rect 13905 12610 13971 12613
rect 15840 12610 16000 12640
rect 13905 12608 16000 12610
rect 13905 12552 13910 12608
rect 13966 12552 16000 12608
rect 13905 12550 16000 12552
rect 13905 12547 13971 12550
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 15840 12520 16000 12550
rect 12940 12479 13256 12480
rect 0 12338 160 12368
rect 841 12338 907 12341
rect 0 12336 907 12338
rect 0 12280 846 12336
rect 902 12280 907 12336
rect 0 12278 907 12280
rect 0 12248 160 12278
rect 841 12275 907 12278
rect 11789 12338 11855 12341
rect 15840 12338 16000 12368
rect 11789 12336 16000 12338
rect 11789 12280 11794 12336
rect 11850 12280 16000 12336
rect 11789 12278 16000 12280
rect 11789 12275 11855 12278
rect 15840 12248 16000 12278
rect 7741 12202 7807 12205
rect 13261 12202 13327 12205
rect 14038 12202 14044 12204
rect 7741 12200 12450 12202
rect 7741 12144 7746 12200
rect 7802 12144 12450 12200
rect 7741 12142 12450 12144
rect 7741 12139 7807 12142
rect 12390 12066 12450 12142
rect 13261 12200 14044 12202
rect 13261 12144 13266 12200
rect 13322 12144 14044 12200
rect 13261 12142 14044 12144
rect 13261 12139 13327 12142
rect 14038 12140 14044 12142
rect 14108 12140 14114 12204
rect 14273 12066 14339 12069
rect 12390 12064 14339 12066
rect 12390 12008 14278 12064
rect 14334 12008 14339 12064
rect 12390 12006 14339 12008
rect 14273 12003 14339 12006
rect 15101 12066 15167 12069
rect 15840 12066 16000 12096
rect 15101 12064 16000 12066
rect 15101 12008 15106 12064
rect 15162 12008 16000 12064
rect 15101 12006 16000 12008
rect 15101 12003 15167 12006
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 15840 11976 16000 12006
rect 14653 11935 14969 11936
rect 13721 11932 13787 11933
rect 13670 11868 13676 11932
rect 13740 11930 13787 11932
rect 13740 11928 13832 11930
rect 13782 11872 13832 11928
rect 13740 11870 13832 11872
rect 13740 11868 13787 11870
rect 13721 11867 13787 11868
rect 13486 11732 13492 11796
rect 13556 11794 13562 11796
rect 13905 11794 13971 11797
rect 13556 11792 13971 11794
rect 13556 11736 13910 11792
rect 13966 11736 13971 11792
rect 13556 11734 13971 11736
rect 13556 11732 13562 11734
rect 13905 11731 13971 11734
rect 14181 11794 14247 11797
rect 15840 11794 16000 11824
rect 14181 11792 16000 11794
rect 14181 11736 14186 11792
rect 14242 11736 16000 11792
rect 14181 11734 16000 11736
rect 14181 11731 14247 11734
rect 15840 11704 16000 11734
rect 7465 11658 7531 11661
rect 8845 11658 8911 11661
rect 7465 11656 8911 11658
rect 7465 11600 7470 11656
rect 7526 11600 8850 11656
rect 8906 11600 8911 11656
rect 7465 11598 8911 11600
rect 7465 11595 7531 11598
rect 8845 11595 8911 11598
rect 0 11522 160 11552
rect 841 11522 907 11525
rect 0 11520 907 11522
rect 0 11464 846 11520
rect 902 11464 907 11520
rect 0 11462 907 11464
rect 0 11432 160 11462
rect 841 11459 907 11462
rect 14641 11522 14707 11525
rect 15840 11522 16000 11552
rect 14641 11520 16000 11522
rect 14641 11464 14646 11520
rect 14702 11464 16000 11520
rect 14641 11462 16000 11464
rect 14641 11459 14707 11462
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 15840 11432 16000 11462
rect 12940 11391 13256 11392
rect 11881 11250 11947 11253
rect 15840 11250 16000 11280
rect 11881 11248 16000 11250
rect 11881 11192 11886 11248
rect 11942 11192 16000 11248
rect 11881 11190 16000 11192
rect 11881 11187 11947 11190
rect 15840 11160 16000 11190
rect 14460 11054 15210 11114
rect 1577 10978 1643 10981
rect 798 10976 1643 10978
rect 798 10920 1582 10976
rect 1638 10920 1643 10976
rect 798 10918 1643 10920
rect 0 10706 160 10736
rect 798 10706 858 10918
rect 1577 10915 1643 10918
rect 11697 10978 11763 10981
rect 14460 10978 14520 11054
rect 11697 10976 14520 10978
rect 11697 10920 11702 10976
rect 11758 10920 14520 10976
rect 11697 10918 14520 10920
rect 15150 10978 15210 11054
rect 15840 10978 16000 11008
rect 15150 10918 16000 10978
rect 11697 10915 11763 10918
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 15840 10888 16000 10918
rect 14653 10847 14969 10848
rect 0 10646 858 10706
rect 0 10616 160 10646
rect 2262 10644 2268 10708
rect 2332 10706 2338 10708
rect 8845 10706 8911 10709
rect 2332 10704 8911 10706
rect 2332 10648 8850 10704
rect 8906 10648 8911 10704
rect 2332 10646 8911 10648
rect 2332 10644 2338 10646
rect 8845 10643 8911 10646
rect 11053 10706 11119 10709
rect 15840 10706 16000 10736
rect 11053 10704 16000 10706
rect 11053 10648 11058 10704
rect 11114 10648 16000 10704
rect 11053 10646 16000 10648
rect 11053 10643 11119 10646
rect 15840 10616 16000 10646
rect 6821 10570 6887 10573
rect 8477 10570 8543 10573
rect 6821 10568 8543 10570
rect 6821 10512 6826 10568
rect 6882 10512 8482 10568
rect 8538 10512 8543 10568
rect 6821 10510 8543 10512
rect 6821 10507 6887 10510
rect 8477 10507 8543 10510
rect 10317 10570 10383 10573
rect 13629 10570 13695 10573
rect 10317 10568 13695 10570
rect 10317 10512 10322 10568
rect 10378 10512 13634 10568
rect 13690 10512 13695 10568
rect 10317 10510 13695 10512
rect 10317 10507 10383 10510
rect 13629 10507 13695 10510
rect 14181 10434 14247 10437
rect 15840 10434 16000 10464
rect 14181 10432 16000 10434
rect 14181 10376 14186 10432
rect 14242 10376 16000 10432
rect 14181 10374 16000 10376
rect 14181 10371 14247 10374
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 15840 10344 16000 10374
rect 12940 10303 13256 10304
rect 12709 10162 12775 10165
rect 13905 10162 13971 10165
rect 12709 10160 13971 10162
rect 12709 10104 12714 10160
rect 12770 10104 13910 10160
rect 13966 10104 13971 10160
rect 12709 10102 13971 10104
rect 12709 10099 12775 10102
rect 13905 10099 13971 10102
rect 15101 10162 15167 10165
rect 15840 10162 16000 10192
rect 15101 10160 16000 10162
rect 15101 10104 15106 10160
rect 15162 10104 16000 10160
rect 15101 10102 16000 10104
rect 15101 10099 15167 10102
rect 15840 10072 16000 10102
rect 10593 10026 10659 10029
rect 12801 10028 12867 10029
rect 12750 10026 12756 10028
rect 10593 10024 12450 10026
rect 10593 9968 10598 10024
rect 10654 9968 12450 10024
rect 10593 9966 12450 9968
rect 12710 9966 12756 10026
rect 12820 10024 12867 10028
rect 12862 9968 12867 10024
rect 10593 9963 10659 9966
rect 0 9890 160 9920
rect 1025 9890 1091 9893
rect 0 9888 1091 9890
rect 0 9832 1030 9888
rect 1086 9832 1091 9888
rect 0 9830 1091 9832
rect 0 9800 160 9830
rect 1025 9827 1091 9830
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 11646 9692 11652 9756
rect 11716 9754 11722 9756
rect 12249 9754 12315 9757
rect 11716 9752 12315 9754
rect 11716 9696 12254 9752
rect 12310 9696 12315 9752
rect 11716 9694 12315 9696
rect 11716 9692 11722 9694
rect 12249 9691 12315 9694
rect 1577 9618 1643 9621
rect 1761 9620 1827 9621
rect 62 9616 1643 9618
rect 62 9560 1582 9616
rect 1638 9560 1643 9616
rect 62 9558 1643 9560
rect 62 9346 122 9558
rect 1577 9555 1643 9558
rect 1710 9556 1716 9620
rect 1780 9618 1827 9620
rect 12157 9618 12223 9621
rect 1780 9616 12223 9618
rect 1822 9560 12162 9616
rect 12218 9560 12223 9616
rect 1780 9558 12223 9560
rect 1780 9556 1827 9558
rect 1761 9555 1827 9556
rect 12157 9555 12223 9558
rect 1853 9482 1919 9485
rect 11881 9482 11947 9485
rect 1853 9480 11947 9482
rect 1853 9424 1858 9480
rect 1914 9424 11886 9480
rect 11942 9424 11947 9480
rect 1853 9422 11947 9424
rect 12390 9482 12450 9966
rect 12750 9964 12756 9966
rect 12820 9964 12867 9968
rect 12801 9963 12867 9964
rect 15469 9890 15535 9893
rect 15840 9890 16000 9920
rect 15469 9888 16000 9890
rect 15469 9832 15474 9888
rect 15530 9832 16000 9888
rect 15469 9830 16000 9832
rect 15469 9827 15535 9830
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 15840 9800 16000 9830
rect 14653 9759 14969 9760
rect 14273 9618 14339 9621
rect 15840 9618 16000 9648
rect 14273 9616 16000 9618
rect 14273 9560 14278 9616
rect 14334 9560 16000 9616
rect 14273 9558 16000 9560
rect 14273 9555 14339 9558
rect 15840 9528 16000 9558
rect 13445 9482 13511 9485
rect 12390 9480 13511 9482
rect 12390 9424 13450 9480
rect 13506 9424 13511 9480
rect 12390 9422 13511 9424
rect 1853 9419 1919 9422
rect 11881 9419 11947 9422
rect 13445 9419 13511 9422
rect 11237 9346 11303 9349
rect 11646 9346 11652 9348
rect 62 9286 306 9346
rect 0 9074 160 9104
rect 246 9074 306 9286
rect 11237 9344 11652 9346
rect 11237 9288 11242 9344
rect 11298 9288 11652 9344
rect 11237 9286 11652 9288
rect 11237 9283 11303 9286
rect 11646 9284 11652 9286
rect 11716 9284 11722 9348
rect 11789 9346 11855 9349
rect 13813 9346 13879 9349
rect 15840 9346 16000 9376
rect 11789 9344 12818 9346
rect 11789 9288 11794 9344
rect 11850 9288 12818 9344
rect 11789 9286 12818 9288
rect 11789 9283 11855 9286
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 10317 9210 10383 9213
rect 11697 9210 11763 9213
rect 10317 9208 11763 9210
rect 10317 9152 10322 9208
rect 10378 9152 11702 9208
rect 11758 9152 11763 9208
rect 10317 9150 11763 9152
rect 10317 9147 10383 9150
rect 11697 9147 11763 9150
rect 12341 9208 12407 9213
rect 12341 9152 12346 9208
rect 12402 9152 12407 9208
rect 12341 9147 12407 9152
rect 0 9014 306 9074
rect 10869 9074 10935 9077
rect 11421 9074 11487 9077
rect 10869 9072 11487 9074
rect 10869 9016 10874 9072
rect 10930 9016 11426 9072
rect 11482 9016 11487 9072
rect 10869 9014 11487 9016
rect 0 8984 160 9014
rect 10869 9011 10935 9014
rect 11421 9011 11487 9014
rect 11973 9074 12039 9077
rect 12198 9074 12204 9076
rect 11973 9072 12204 9074
rect 11973 9016 11978 9072
rect 12034 9016 12204 9072
rect 11973 9014 12204 9016
rect 11973 9011 12039 9014
rect 12198 9012 12204 9014
rect 12268 9012 12274 9076
rect 7097 8938 7163 8941
rect 10133 8938 10199 8941
rect 7097 8936 10199 8938
rect 7097 8880 7102 8936
rect 7158 8880 10138 8936
rect 10194 8880 10199 8936
rect 7097 8878 10199 8880
rect 7097 8875 7163 8878
rect 10133 8875 10199 8878
rect 11145 8938 11211 8941
rect 11973 8938 12039 8941
rect 11145 8936 12039 8938
rect 11145 8880 11150 8936
rect 11206 8880 11978 8936
rect 12034 8880 12039 8936
rect 11145 8878 12039 8880
rect 12344 8938 12404 9147
rect 12758 9074 12818 9286
rect 13813 9344 16000 9346
rect 13813 9288 13818 9344
rect 13874 9288 16000 9344
rect 13813 9286 16000 9288
rect 13813 9283 13879 9286
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 15840 9256 16000 9286
rect 12940 9215 13256 9216
rect 15840 9074 16000 9104
rect 12758 9014 16000 9074
rect 15840 8984 16000 9014
rect 12344 8878 15164 8938
rect 11145 8875 11211 8878
rect 11973 8875 12039 8878
rect 15104 8802 15164 8878
rect 15840 8802 16000 8832
rect 15104 8742 16000 8802
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 15840 8712 16000 8742
rect 14653 8671 14969 8672
rect 12198 8604 12204 8668
rect 12268 8666 12274 8668
rect 12709 8666 12775 8669
rect 12268 8664 12775 8666
rect 12268 8608 12714 8664
rect 12770 8608 12775 8664
rect 12268 8606 12775 8608
rect 12268 8604 12274 8606
rect 12709 8603 12775 8606
rect 7189 8530 7255 8533
rect 9857 8530 9923 8533
rect 7189 8528 9923 8530
rect 7189 8472 7194 8528
rect 7250 8472 9862 8528
rect 9918 8472 9923 8528
rect 7189 8470 9923 8472
rect 7189 8467 7255 8470
rect 9857 8467 9923 8470
rect 11513 8530 11579 8533
rect 15840 8530 16000 8560
rect 11513 8528 16000 8530
rect 11513 8472 11518 8528
rect 11574 8472 16000 8528
rect 11513 8470 16000 8472
rect 11513 8467 11579 8470
rect 15840 8440 16000 8470
rect 5441 8394 5507 8397
rect 12801 8394 12867 8397
rect 5441 8392 12867 8394
rect 5441 8336 5446 8392
rect 5502 8336 12806 8392
rect 12862 8336 12867 8392
rect 5441 8334 12867 8336
rect 5441 8331 5507 8334
rect 12801 8331 12867 8334
rect 0 8258 160 8288
rect 1669 8258 1735 8261
rect 0 8256 1735 8258
rect 0 8200 1674 8256
rect 1730 8200 1735 8256
rect 0 8198 1735 8200
rect 0 8168 160 8198
rect 1669 8195 1735 8198
rect 14273 8258 14339 8261
rect 15840 8258 16000 8288
rect 14273 8256 16000 8258
rect 14273 8200 14278 8256
rect 14334 8200 16000 8256
rect 14273 8198 16000 8200
rect 14273 8195 14339 8198
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 15840 8168 16000 8198
rect 12940 8127 13256 8128
rect 13353 7986 13419 7989
rect 15840 7986 16000 8016
rect 13353 7984 16000 7986
rect 13353 7928 13358 7984
rect 13414 7928 16000 7984
rect 13353 7926 16000 7928
rect 13353 7923 13419 7926
rect 15840 7896 16000 7926
rect 11329 7850 11395 7853
rect 12157 7850 12223 7853
rect 11329 7848 12223 7850
rect 11329 7792 11334 7848
rect 11390 7792 12162 7848
rect 12218 7792 12223 7848
rect 11329 7790 12223 7792
rect 11329 7787 11395 7790
rect 12157 7787 12223 7790
rect 15101 7714 15167 7717
rect 15840 7714 16000 7744
rect 15101 7712 16000 7714
rect 15101 7656 15106 7712
rect 15162 7656 16000 7712
rect 15101 7654 16000 7656
rect 15101 7651 15167 7654
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 15840 7624 16000 7654
rect 14653 7583 14969 7584
rect 0 7442 160 7472
rect 841 7442 907 7445
rect 0 7440 907 7442
rect 0 7384 846 7440
rect 902 7384 907 7440
rect 0 7382 907 7384
rect 0 7352 160 7382
rect 841 7379 907 7382
rect 13721 7442 13787 7445
rect 15840 7442 16000 7472
rect 13721 7440 16000 7442
rect 13721 7384 13726 7440
rect 13782 7384 16000 7440
rect 13721 7382 16000 7384
rect 13721 7379 13787 7382
rect 15840 7352 16000 7382
rect 13721 7170 13787 7173
rect 15840 7170 16000 7200
rect 13721 7168 16000 7170
rect 13721 7112 13726 7168
rect 13782 7112 16000 7168
rect 13721 7110 16000 7112
rect 13721 7107 13787 7110
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 15840 7080 16000 7110
rect 12940 7039 13256 7040
rect 12341 6898 12407 6901
rect 15840 6898 16000 6928
rect 12341 6896 16000 6898
rect 12341 6840 12346 6896
rect 12402 6840 16000 6896
rect 12341 6838 16000 6840
rect 12341 6835 12407 6838
rect 15840 6808 16000 6838
rect 9029 6762 9095 6765
rect 13629 6762 13695 6765
rect 9029 6760 13695 6762
rect 9029 6704 9034 6760
rect 9090 6704 13634 6760
rect 13690 6704 13695 6760
rect 9029 6702 13695 6704
rect 9029 6699 9095 6702
rect 13629 6699 13695 6702
rect 0 6626 160 6656
rect 841 6626 907 6629
rect 0 6624 907 6626
rect 0 6568 846 6624
rect 902 6568 907 6624
rect 0 6566 907 6568
rect 0 6536 160 6566
rect 841 6563 907 6566
rect 15101 6626 15167 6629
rect 15840 6626 16000 6656
rect 15101 6624 16000 6626
rect 15101 6568 15106 6624
rect 15162 6568 16000 6624
rect 15101 6566 16000 6568
rect 15101 6563 15167 6566
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 15840 6536 16000 6566
rect 14653 6495 14969 6496
rect 12433 6354 12499 6357
rect 12893 6354 12959 6357
rect 12433 6352 12959 6354
rect 12433 6296 12438 6352
rect 12494 6296 12898 6352
rect 12954 6296 12959 6352
rect 12433 6294 12959 6296
rect 12433 6291 12499 6294
rect 12893 6291 12959 6294
rect 14733 6354 14799 6357
rect 15840 6354 16000 6384
rect 14733 6352 16000 6354
rect 14733 6296 14738 6352
rect 14794 6296 16000 6352
rect 14733 6294 16000 6296
rect 14733 6291 14799 6294
rect 15840 6264 16000 6294
rect 9673 6218 9739 6221
rect 13905 6218 13971 6221
rect 9673 6216 13971 6218
rect 9673 6160 9678 6216
rect 9734 6160 13910 6216
rect 13966 6160 13971 6216
rect 9673 6158 13971 6160
rect 9673 6155 9739 6158
rect 13905 6155 13971 6158
rect 14181 6082 14247 6085
rect 15840 6082 16000 6112
rect 14181 6080 16000 6082
rect 14181 6024 14186 6080
rect 14242 6024 16000 6080
rect 14181 6022 16000 6024
rect 14181 6019 14247 6022
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 15840 5992 16000 6022
rect 12940 5951 13256 5952
rect 0 5810 160 5840
rect 841 5810 907 5813
rect 0 5808 907 5810
rect 0 5752 846 5808
rect 902 5752 907 5808
rect 0 5750 907 5752
rect 0 5720 160 5750
rect 841 5747 907 5750
rect 8293 5810 8359 5813
rect 13353 5810 13419 5813
rect 15840 5810 16000 5840
rect 8293 5808 13419 5810
rect 8293 5752 8298 5808
rect 8354 5752 13358 5808
rect 13414 5752 13419 5808
rect 8293 5750 13419 5752
rect 8293 5747 8359 5750
rect 13353 5747 13419 5750
rect 14966 5750 16000 5810
rect 2497 5674 2563 5677
rect 13905 5674 13971 5677
rect 2497 5672 13971 5674
rect 2497 5616 2502 5672
rect 2558 5616 13910 5672
rect 13966 5616 13971 5672
rect 2497 5614 13971 5616
rect 2497 5611 2563 5614
rect 13905 5611 13971 5614
rect 14181 5674 14247 5677
rect 14966 5674 15026 5750
rect 15840 5720 16000 5750
rect 14181 5672 15026 5674
rect 14181 5616 14186 5672
rect 14242 5616 15026 5672
rect 14181 5614 15026 5616
rect 14181 5611 14247 5614
rect 15101 5538 15167 5541
rect 15840 5538 16000 5568
rect 15101 5536 16000 5538
rect 15101 5480 15106 5536
rect 15162 5480 16000 5536
rect 15101 5478 16000 5480
rect 15101 5475 15167 5478
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 15840 5448 16000 5478
rect 14653 5407 14969 5408
rect 13721 5266 13787 5269
rect 15840 5266 16000 5296
rect 13721 5264 16000 5266
rect 13721 5208 13726 5264
rect 13782 5208 16000 5264
rect 13721 5206 16000 5208
rect 13721 5203 13787 5206
rect 15840 5176 16000 5206
rect 0 4994 160 5024
rect 841 4994 907 4997
rect 0 4992 907 4994
rect 0 4936 846 4992
rect 902 4936 907 4992
rect 0 4934 907 4936
rect 0 4904 160 4934
rect 841 4931 907 4934
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 0 4178 160 4208
rect 749 4178 815 4181
rect 0 4176 815 4178
rect 0 4120 754 4176
rect 810 4120 815 4176
rect 0 4118 815 4120
rect 0 4088 160 4118
rect 749 4115 815 4118
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 6678 3436 6684 3500
rect 6748 3498 6754 3500
rect 12433 3498 12499 3501
rect 6748 3496 12499 3498
rect 6748 3440 12438 3496
rect 12494 3440 12499 3496
rect 6748 3438 12499 3440
rect 6748 3436 6754 3438
rect 12433 3435 12499 3438
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 10910 2620 10916 2684
rect 10980 2682 10986 2684
rect 11053 2682 11119 2685
rect 11789 2684 11855 2685
rect 11789 2682 11836 2684
rect 10980 2680 11119 2682
rect 10980 2624 11058 2680
rect 11114 2624 11119 2680
rect 10980 2622 11119 2624
rect 11744 2680 11836 2682
rect 11744 2624 11794 2680
rect 11744 2622 11836 2624
rect 10980 2620 10986 2622
rect 11053 2619 11119 2622
rect 11789 2620 11836 2622
rect 11900 2620 11906 2684
rect 11789 2619 11855 2620
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
rect 2659 1664 2975 1665
rect 2659 1600 2665 1664
rect 2729 1600 2745 1664
rect 2809 1600 2825 1664
rect 2889 1600 2905 1664
rect 2969 1600 2975 1664
rect 2659 1599 2975 1600
rect 6086 1664 6402 1665
rect 6086 1600 6092 1664
rect 6156 1600 6172 1664
rect 6236 1600 6252 1664
rect 6316 1600 6332 1664
rect 6396 1600 6402 1664
rect 6086 1599 6402 1600
rect 9513 1664 9829 1665
rect 9513 1600 9519 1664
rect 9583 1600 9599 1664
rect 9663 1600 9679 1664
rect 9743 1600 9759 1664
rect 9823 1600 9829 1664
rect 9513 1599 9829 1600
rect 12940 1664 13256 1665
rect 12940 1600 12946 1664
rect 13010 1600 13026 1664
rect 13090 1600 13106 1664
rect 13170 1600 13186 1664
rect 13250 1600 13256 1664
rect 12940 1599 13256 1600
rect 4613 1322 4679 1325
rect 5349 1324 5415 1325
rect 4838 1322 4844 1324
rect 4613 1320 4844 1322
rect 4613 1264 4618 1320
rect 4674 1264 4844 1320
rect 4613 1262 4844 1264
rect 4613 1259 4679 1262
rect 4838 1260 4844 1262
rect 4908 1260 4914 1324
rect 5349 1322 5396 1324
rect 5304 1320 5396 1322
rect 5304 1264 5354 1320
rect 5304 1262 5396 1264
rect 5349 1260 5396 1262
rect 5460 1260 5466 1324
rect 5349 1259 5415 1260
rect 4372 1120 4688 1121
rect 4372 1056 4378 1120
rect 4442 1056 4458 1120
rect 4522 1056 4538 1120
rect 4602 1056 4618 1120
rect 4682 1056 4688 1120
rect 4372 1055 4688 1056
rect 7799 1120 8115 1121
rect 7799 1056 7805 1120
rect 7869 1056 7885 1120
rect 7949 1056 7965 1120
rect 8029 1056 8045 1120
rect 8109 1056 8115 1120
rect 7799 1055 8115 1056
rect 11226 1120 11542 1121
rect 11226 1056 11232 1120
rect 11296 1056 11312 1120
rect 11376 1056 11392 1120
rect 11456 1056 11472 1120
rect 11536 1056 11542 1120
rect 11226 1055 11542 1056
rect 14653 1120 14969 1121
rect 14653 1056 14659 1120
rect 14723 1056 14739 1120
rect 14803 1056 14819 1120
rect 14883 1056 14899 1120
rect 14963 1056 14969 1120
rect 14653 1055 14969 1056
<< via3 >>
rect 4378 43548 4442 43552
rect 4378 43492 4382 43548
rect 4382 43492 4438 43548
rect 4438 43492 4442 43548
rect 4378 43488 4442 43492
rect 4458 43548 4522 43552
rect 4458 43492 4462 43548
rect 4462 43492 4518 43548
rect 4518 43492 4522 43548
rect 4458 43488 4522 43492
rect 4538 43548 4602 43552
rect 4538 43492 4542 43548
rect 4542 43492 4598 43548
rect 4598 43492 4602 43548
rect 4538 43488 4602 43492
rect 4618 43548 4682 43552
rect 4618 43492 4622 43548
rect 4622 43492 4678 43548
rect 4678 43492 4682 43548
rect 4618 43488 4682 43492
rect 7805 43548 7869 43552
rect 7805 43492 7809 43548
rect 7809 43492 7865 43548
rect 7865 43492 7869 43548
rect 7805 43488 7869 43492
rect 7885 43548 7949 43552
rect 7885 43492 7889 43548
rect 7889 43492 7945 43548
rect 7945 43492 7949 43548
rect 7885 43488 7949 43492
rect 7965 43548 8029 43552
rect 7965 43492 7969 43548
rect 7969 43492 8025 43548
rect 8025 43492 8029 43548
rect 7965 43488 8029 43492
rect 8045 43548 8109 43552
rect 8045 43492 8049 43548
rect 8049 43492 8105 43548
rect 8105 43492 8109 43548
rect 8045 43488 8109 43492
rect 11232 43548 11296 43552
rect 11232 43492 11236 43548
rect 11236 43492 11292 43548
rect 11292 43492 11296 43548
rect 11232 43488 11296 43492
rect 11312 43548 11376 43552
rect 11312 43492 11316 43548
rect 11316 43492 11372 43548
rect 11372 43492 11376 43548
rect 11312 43488 11376 43492
rect 11392 43548 11456 43552
rect 11392 43492 11396 43548
rect 11396 43492 11452 43548
rect 11452 43492 11456 43548
rect 11392 43488 11456 43492
rect 11472 43548 11536 43552
rect 11472 43492 11476 43548
rect 11476 43492 11532 43548
rect 11532 43492 11536 43548
rect 11472 43488 11536 43492
rect 14659 43548 14723 43552
rect 14659 43492 14663 43548
rect 14663 43492 14719 43548
rect 14719 43492 14723 43548
rect 14659 43488 14723 43492
rect 14739 43548 14803 43552
rect 14739 43492 14743 43548
rect 14743 43492 14799 43548
rect 14799 43492 14803 43548
rect 14739 43488 14803 43492
rect 14819 43548 14883 43552
rect 14819 43492 14823 43548
rect 14823 43492 14879 43548
rect 14879 43492 14883 43548
rect 14819 43488 14883 43492
rect 14899 43548 14963 43552
rect 14899 43492 14903 43548
rect 14903 43492 14959 43548
rect 14959 43492 14963 43548
rect 14899 43488 14963 43492
rect 2665 43004 2729 43008
rect 2665 42948 2669 43004
rect 2669 42948 2725 43004
rect 2725 42948 2729 43004
rect 2665 42944 2729 42948
rect 2745 43004 2809 43008
rect 2745 42948 2749 43004
rect 2749 42948 2805 43004
rect 2805 42948 2809 43004
rect 2745 42944 2809 42948
rect 2825 43004 2889 43008
rect 2825 42948 2829 43004
rect 2829 42948 2885 43004
rect 2885 42948 2889 43004
rect 2825 42944 2889 42948
rect 2905 43004 2969 43008
rect 2905 42948 2909 43004
rect 2909 42948 2965 43004
rect 2965 42948 2969 43004
rect 2905 42944 2969 42948
rect 6092 43004 6156 43008
rect 6092 42948 6096 43004
rect 6096 42948 6152 43004
rect 6152 42948 6156 43004
rect 6092 42944 6156 42948
rect 6172 43004 6236 43008
rect 6172 42948 6176 43004
rect 6176 42948 6232 43004
rect 6232 42948 6236 43004
rect 6172 42944 6236 42948
rect 6252 43004 6316 43008
rect 6252 42948 6256 43004
rect 6256 42948 6312 43004
rect 6312 42948 6316 43004
rect 6252 42944 6316 42948
rect 6332 43004 6396 43008
rect 6332 42948 6336 43004
rect 6336 42948 6392 43004
rect 6392 42948 6396 43004
rect 6332 42944 6396 42948
rect 9519 43004 9583 43008
rect 9519 42948 9523 43004
rect 9523 42948 9579 43004
rect 9579 42948 9583 43004
rect 9519 42944 9583 42948
rect 9599 43004 9663 43008
rect 9599 42948 9603 43004
rect 9603 42948 9659 43004
rect 9659 42948 9663 43004
rect 9599 42944 9663 42948
rect 9679 43004 9743 43008
rect 9679 42948 9683 43004
rect 9683 42948 9739 43004
rect 9739 42948 9743 43004
rect 9679 42944 9743 42948
rect 9759 43004 9823 43008
rect 9759 42948 9763 43004
rect 9763 42948 9819 43004
rect 9819 42948 9823 43004
rect 9759 42944 9823 42948
rect 12946 43004 13010 43008
rect 12946 42948 12950 43004
rect 12950 42948 13006 43004
rect 13006 42948 13010 43004
rect 12946 42944 13010 42948
rect 13026 43004 13090 43008
rect 13026 42948 13030 43004
rect 13030 42948 13086 43004
rect 13086 42948 13090 43004
rect 13026 42944 13090 42948
rect 13106 43004 13170 43008
rect 13106 42948 13110 43004
rect 13110 42948 13166 43004
rect 13166 42948 13170 43004
rect 13106 42944 13170 42948
rect 13186 43004 13250 43008
rect 13186 42948 13190 43004
rect 13190 42948 13246 43004
rect 13246 42948 13250 43004
rect 13186 42944 13250 42948
rect 6684 42604 6748 42668
rect 4378 42460 4442 42464
rect 4378 42404 4382 42460
rect 4382 42404 4438 42460
rect 4438 42404 4442 42460
rect 4378 42400 4442 42404
rect 4458 42460 4522 42464
rect 4458 42404 4462 42460
rect 4462 42404 4518 42460
rect 4518 42404 4522 42460
rect 4458 42400 4522 42404
rect 4538 42460 4602 42464
rect 4538 42404 4542 42460
rect 4542 42404 4598 42460
rect 4598 42404 4602 42460
rect 4538 42400 4602 42404
rect 4618 42460 4682 42464
rect 4618 42404 4622 42460
rect 4622 42404 4678 42460
rect 4678 42404 4682 42460
rect 4618 42400 4682 42404
rect 7805 42460 7869 42464
rect 7805 42404 7809 42460
rect 7809 42404 7865 42460
rect 7865 42404 7869 42460
rect 7805 42400 7869 42404
rect 7885 42460 7949 42464
rect 7885 42404 7889 42460
rect 7889 42404 7945 42460
rect 7945 42404 7949 42460
rect 7885 42400 7949 42404
rect 7965 42460 8029 42464
rect 7965 42404 7969 42460
rect 7969 42404 8025 42460
rect 8025 42404 8029 42460
rect 7965 42400 8029 42404
rect 8045 42460 8109 42464
rect 8045 42404 8049 42460
rect 8049 42404 8105 42460
rect 8105 42404 8109 42460
rect 8045 42400 8109 42404
rect 11232 42460 11296 42464
rect 11232 42404 11236 42460
rect 11236 42404 11292 42460
rect 11292 42404 11296 42460
rect 11232 42400 11296 42404
rect 11312 42460 11376 42464
rect 11312 42404 11316 42460
rect 11316 42404 11372 42460
rect 11372 42404 11376 42460
rect 11312 42400 11376 42404
rect 11392 42460 11456 42464
rect 11392 42404 11396 42460
rect 11396 42404 11452 42460
rect 11452 42404 11456 42460
rect 11392 42400 11456 42404
rect 11472 42460 11536 42464
rect 11472 42404 11476 42460
rect 11476 42404 11532 42460
rect 11532 42404 11536 42460
rect 11472 42400 11536 42404
rect 14659 42460 14723 42464
rect 14659 42404 14663 42460
rect 14663 42404 14719 42460
rect 14719 42404 14723 42460
rect 14659 42400 14723 42404
rect 14739 42460 14803 42464
rect 14739 42404 14743 42460
rect 14743 42404 14799 42460
rect 14799 42404 14803 42460
rect 14739 42400 14803 42404
rect 14819 42460 14883 42464
rect 14819 42404 14823 42460
rect 14823 42404 14879 42460
rect 14879 42404 14883 42460
rect 14819 42400 14883 42404
rect 14899 42460 14963 42464
rect 14899 42404 14903 42460
rect 14903 42404 14959 42460
rect 14959 42404 14963 42460
rect 14899 42400 14963 42404
rect 2665 41916 2729 41920
rect 2665 41860 2669 41916
rect 2669 41860 2725 41916
rect 2725 41860 2729 41916
rect 2665 41856 2729 41860
rect 2745 41916 2809 41920
rect 2745 41860 2749 41916
rect 2749 41860 2805 41916
rect 2805 41860 2809 41916
rect 2745 41856 2809 41860
rect 2825 41916 2889 41920
rect 2825 41860 2829 41916
rect 2829 41860 2885 41916
rect 2885 41860 2889 41916
rect 2825 41856 2889 41860
rect 2905 41916 2969 41920
rect 2905 41860 2909 41916
rect 2909 41860 2965 41916
rect 2965 41860 2969 41916
rect 2905 41856 2969 41860
rect 6092 41916 6156 41920
rect 6092 41860 6096 41916
rect 6096 41860 6152 41916
rect 6152 41860 6156 41916
rect 6092 41856 6156 41860
rect 6172 41916 6236 41920
rect 6172 41860 6176 41916
rect 6176 41860 6232 41916
rect 6232 41860 6236 41916
rect 6172 41856 6236 41860
rect 6252 41916 6316 41920
rect 6252 41860 6256 41916
rect 6256 41860 6312 41916
rect 6312 41860 6316 41916
rect 6252 41856 6316 41860
rect 6332 41916 6396 41920
rect 6332 41860 6336 41916
rect 6336 41860 6392 41916
rect 6392 41860 6396 41916
rect 6332 41856 6396 41860
rect 9519 41916 9583 41920
rect 9519 41860 9523 41916
rect 9523 41860 9579 41916
rect 9579 41860 9583 41916
rect 9519 41856 9583 41860
rect 9599 41916 9663 41920
rect 9599 41860 9603 41916
rect 9603 41860 9659 41916
rect 9659 41860 9663 41916
rect 9599 41856 9663 41860
rect 9679 41916 9743 41920
rect 9679 41860 9683 41916
rect 9683 41860 9739 41916
rect 9739 41860 9743 41916
rect 9679 41856 9743 41860
rect 9759 41916 9823 41920
rect 9759 41860 9763 41916
rect 9763 41860 9819 41916
rect 9819 41860 9823 41916
rect 9759 41856 9823 41860
rect 12946 41916 13010 41920
rect 12946 41860 12950 41916
rect 12950 41860 13006 41916
rect 13006 41860 13010 41916
rect 12946 41856 13010 41860
rect 13026 41916 13090 41920
rect 13026 41860 13030 41916
rect 13030 41860 13086 41916
rect 13086 41860 13090 41916
rect 13026 41856 13090 41860
rect 13106 41916 13170 41920
rect 13106 41860 13110 41916
rect 13110 41860 13166 41916
rect 13166 41860 13170 41916
rect 13106 41856 13170 41860
rect 13186 41916 13250 41920
rect 13186 41860 13190 41916
rect 13190 41860 13246 41916
rect 13246 41860 13250 41916
rect 13186 41856 13250 41860
rect 2268 41652 2332 41716
rect 4844 41516 4908 41580
rect 7420 41516 7484 41580
rect 5396 41380 5460 41444
rect 10916 41440 10980 41444
rect 10916 41384 10966 41440
rect 10966 41384 10980 41440
rect 10916 41380 10980 41384
rect 4378 41372 4442 41376
rect 4378 41316 4382 41372
rect 4382 41316 4438 41372
rect 4438 41316 4442 41372
rect 4378 41312 4442 41316
rect 4458 41372 4522 41376
rect 4458 41316 4462 41372
rect 4462 41316 4518 41372
rect 4518 41316 4522 41372
rect 4458 41312 4522 41316
rect 4538 41372 4602 41376
rect 4538 41316 4542 41372
rect 4542 41316 4598 41372
rect 4598 41316 4602 41372
rect 4538 41312 4602 41316
rect 4618 41372 4682 41376
rect 4618 41316 4622 41372
rect 4622 41316 4678 41372
rect 4678 41316 4682 41372
rect 4618 41312 4682 41316
rect 7805 41372 7869 41376
rect 7805 41316 7809 41372
rect 7809 41316 7865 41372
rect 7865 41316 7869 41372
rect 7805 41312 7869 41316
rect 7885 41372 7949 41376
rect 7885 41316 7889 41372
rect 7889 41316 7945 41372
rect 7945 41316 7949 41372
rect 7885 41312 7949 41316
rect 7965 41372 8029 41376
rect 7965 41316 7969 41372
rect 7969 41316 8025 41372
rect 8025 41316 8029 41372
rect 7965 41312 8029 41316
rect 8045 41372 8109 41376
rect 8045 41316 8049 41372
rect 8049 41316 8105 41372
rect 8105 41316 8109 41372
rect 8045 41312 8109 41316
rect 11232 41372 11296 41376
rect 11232 41316 11236 41372
rect 11236 41316 11292 41372
rect 11292 41316 11296 41372
rect 11232 41312 11296 41316
rect 11312 41372 11376 41376
rect 11312 41316 11316 41372
rect 11316 41316 11372 41372
rect 11372 41316 11376 41372
rect 11312 41312 11376 41316
rect 11392 41372 11456 41376
rect 11392 41316 11396 41372
rect 11396 41316 11452 41372
rect 11452 41316 11456 41372
rect 11392 41312 11456 41316
rect 11472 41372 11536 41376
rect 11472 41316 11476 41372
rect 11476 41316 11532 41372
rect 11532 41316 11536 41372
rect 11472 41312 11536 41316
rect 14659 41372 14723 41376
rect 14659 41316 14663 41372
rect 14663 41316 14719 41372
rect 14719 41316 14723 41372
rect 14659 41312 14723 41316
rect 14739 41372 14803 41376
rect 14739 41316 14743 41372
rect 14743 41316 14799 41372
rect 14799 41316 14803 41372
rect 14739 41312 14803 41316
rect 14819 41372 14883 41376
rect 14819 41316 14823 41372
rect 14823 41316 14879 41372
rect 14879 41316 14883 41372
rect 14819 41312 14883 41316
rect 14899 41372 14963 41376
rect 14899 41316 14903 41372
rect 14903 41316 14959 41372
rect 14959 41316 14963 41372
rect 14899 41312 14963 41316
rect 2665 40828 2729 40832
rect 2665 40772 2669 40828
rect 2669 40772 2725 40828
rect 2725 40772 2729 40828
rect 2665 40768 2729 40772
rect 2745 40828 2809 40832
rect 2745 40772 2749 40828
rect 2749 40772 2805 40828
rect 2805 40772 2809 40828
rect 2745 40768 2809 40772
rect 2825 40828 2889 40832
rect 2825 40772 2829 40828
rect 2829 40772 2885 40828
rect 2885 40772 2889 40828
rect 2825 40768 2889 40772
rect 2905 40828 2969 40832
rect 2905 40772 2909 40828
rect 2909 40772 2965 40828
rect 2965 40772 2969 40828
rect 2905 40768 2969 40772
rect 6092 40828 6156 40832
rect 6092 40772 6096 40828
rect 6096 40772 6152 40828
rect 6152 40772 6156 40828
rect 6092 40768 6156 40772
rect 6172 40828 6236 40832
rect 6172 40772 6176 40828
rect 6176 40772 6232 40828
rect 6232 40772 6236 40828
rect 6172 40768 6236 40772
rect 6252 40828 6316 40832
rect 6252 40772 6256 40828
rect 6256 40772 6312 40828
rect 6312 40772 6316 40828
rect 6252 40768 6316 40772
rect 6332 40828 6396 40832
rect 6332 40772 6336 40828
rect 6336 40772 6392 40828
rect 6392 40772 6396 40828
rect 6332 40768 6396 40772
rect 9519 40828 9583 40832
rect 9519 40772 9523 40828
rect 9523 40772 9579 40828
rect 9579 40772 9583 40828
rect 9519 40768 9583 40772
rect 9599 40828 9663 40832
rect 9599 40772 9603 40828
rect 9603 40772 9659 40828
rect 9659 40772 9663 40828
rect 9599 40768 9663 40772
rect 9679 40828 9743 40832
rect 9679 40772 9683 40828
rect 9683 40772 9739 40828
rect 9739 40772 9743 40828
rect 9679 40768 9743 40772
rect 9759 40828 9823 40832
rect 9759 40772 9763 40828
rect 9763 40772 9819 40828
rect 9819 40772 9823 40828
rect 9759 40768 9823 40772
rect 12946 40828 13010 40832
rect 12946 40772 12950 40828
rect 12950 40772 13006 40828
rect 13006 40772 13010 40828
rect 12946 40768 13010 40772
rect 13026 40828 13090 40832
rect 13026 40772 13030 40828
rect 13030 40772 13086 40828
rect 13086 40772 13090 40828
rect 13026 40768 13090 40772
rect 13106 40828 13170 40832
rect 13106 40772 13110 40828
rect 13110 40772 13166 40828
rect 13166 40772 13170 40828
rect 13106 40768 13170 40772
rect 13186 40828 13250 40832
rect 13186 40772 13190 40828
rect 13190 40772 13246 40828
rect 13246 40772 13250 40828
rect 13186 40768 13250 40772
rect 4378 40284 4442 40288
rect 4378 40228 4382 40284
rect 4382 40228 4438 40284
rect 4438 40228 4442 40284
rect 4378 40224 4442 40228
rect 4458 40284 4522 40288
rect 4458 40228 4462 40284
rect 4462 40228 4518 40284
rect 4518 40228 4522 40284
rect 4458 40224 4522 40228
rect 4538 40284 4602 40288
rect 4538 40228 4542 40284
rect 4542 40228 4598 40284
rect 4598 40228 4602 40284
rect 4538 40224 4602 40228
rect 4618 40284 4682 40288
rect 4618 40228 4622 40284
rect 4622 40228 4678 40284
rect 4678 40228 4682 40284
rect 4618 40224 4682 40228
rect 7805 40284 7869 40288
rect 7805 40228 7809 40284
rect 7809 40228 7865 40284
rect 7865 40228 7869 40284
rect 7805 40224 7869 40228
rect 7885 40284 7949 40288
rect 7885 40228 7889 40284
rect 7889 40228 7945 40284
rect 7945 40228 7949 40284
rect 7885 40224 7949 40228
rect 7965 40284 8029 40288
rect 7965 40228 7969 40284
rect 7969 40228 8025 40284
rect 8025 40228 8029 40284
rect 7965 40224 8029 40228
rect 8045 40284 8109 40288
rect 8045 40228 8049 40284
rect 8049 40228 8105 40284
rect 8105 40228 8109 40284
rect 8045 40224 8109 40228
rect 11232 40284 11296 40288
rect 11232 40228 11236 40284
rect 11236 40228 11292 40284
rect 11292 40228 11296 40284
rect 11232 40224 11296 40228
rect 11312 40284 11376 40288
rect 11312 40228 11316 40284
rect 11316 40228 11372 40284
rect 11372 40228 11376 40284
rect 11312 40224 11376 40228
rect 11392 40284 11456 40288
rect 11392 40228 11396 40284
rect 11396 40228 11452 40284
rect 11452 40228 11456 40284
rect 11392 40224 11456 40228
rect 11472 40284 11536 40288
rect 11472 40228 11476 40284
rect 11476 40228 11532 40284
rect 11532 40228 11536 40284
rect 11472 40224 11536 40228
rect 14659 40284 14723 40288
rect 14659 40228 14663 40284
rect 14663 40228 14719 40284
rect 14719 40228 14723 40284
rect 14659 40224 14723 40228
rect 14739 40284 14803 40288
rect 14739 40228 14743 40284
rect 14743 40228 14799 40284
rect 14799 40228 14803 40284
rect 14739 40224 14803 40228
rect 14819 40284 14883 40288
rect 14819 40228 14823 40284
rect 14823 40228 14879 40284
rect 14879 40228 14883 40284
rect 14819 40224 14883 40228
rect 14899 40284 14963 40288
rect 14899 40228 14903 40284
rect 14903 40228 14959 40284
rect 14959 40228 14963 40284
rect 14899 40224 14963 40228
rect 9260 40080 9324 40084
rect 9260 40024 9310 40080
rect 9310 40024 9324 40080
rect 9260 40020 9324 40024
rect 2665 39740 2729 39744
rect 2665 39684 2669 39740
rect 2669 39684 2725 39740
rect 2725 39684 2729 39740
rect 2665 39680 2729 39684
rect 2745 39740 2809 39744
rect 2745 39684 2749 39740
rect 2749 39684 2805 39740
rect 2805 39684 2809 39740
rect 2745 39680 2809 39684
rect 2825 39740 2889 39744
rect 2825 39684 2829 39740
rect 2829 39684 2885 39740
rect 2885 39684 2889 39740
rect 2825 39680 2889 39684
rect 2905 39740 2969 39744
rect 2905 39684 2909 39740
rect 2909 39684 2965 39740
rect 2965 39684 2969 39740
rect 2905 39680 2969 39684
rect 6092 39740 6156 39744
rect 6092 39684 6096 39740
rect 6096 39684 6152 39740
rect 6152 39684 6156 39740
rect 6092 39680 6156 39684
rect 6172 39740 6236 39744
rect 6172 39684 6176 39740
rect 6176 39684 6232 39740
rect 6232 39684 6236 39740
rect 6172 39680 6236 39684
rect 6252 39740 6316 39744
rect 6252 39684 6256 39740
rect 6256 39684 6312 39740
rect 6312 39684 6316 39740
rect 6252 39680 6316 39684
rect 6332 39740 6396 39744
rect 6332 39684 6336 39740
rect 6336 39684 6392 39740
rect 6392 39684 6396 39740
rect 6332 39680 6396 39684
rect 9519 39740 9583 39744
rect 9519 39684 9523 39740
rect 9523 39684 9579 39740
rect 9579 39684 9583 39740
rect 9519 39680 9583 39684
rect 9599 39740 9663 39744
rect 9599 39684 9603 39740
rect 9603 39684 9659 39740
rect 9659 39684 9663 39740
rect 9599 39680 9663 39684
rect 9679 39740 9743 39744
rect 9679 39684 9683 39740
rect 9683 39684 9739 39740
rect 9739 39684 9743 39740
rect 9679 39680 9743 39684
rect 9759 39740 9823 39744
rect 9759 39684 9763 39740
rect 9763 39684 9819 39740
rect 9819 39684 9823 39740
rect 9759 39680 9823 39684
rect 12946 39740 13010 39744
rect 12946 39684 12950 39740
rect 12950 39684 13006 39740
rect 13006 39684 13010 39740
rect 12946 39680 13010 39684
rect 13026 39740 13090 39744
rect 13026 39684 13030 39740
rect 13030 39684 13086 39740
rect 13086 39684 13090 39740
rect 13026 39680 13090 39684
rect 13106 39740 13170 39744
rect 13106 39684 13110 39740
rect 13110 39684 13166 39740
rect 13166 39684 13170 39740
rect 13106 39680 13170 39684
rect 13186 39740 13250 39744
rect 13186 39684 13190 39740
rect 13190 39684 13246 39740
rect 13246 39684 13250 39740
rect 13186 39680 13250 39684
rect 4378 39196 4442 39200
rect 4378 39140 4382 39196
rect 4382 39140 4438 39196
rect 4438 39140 4442 39196
rect 4378 39136 4442 39140
rect 4458 39196 4522 39200
rect 4458 39140 4462 39196
rect 4462 39140 4518 39196
rect 4518 39140 4522 39196
rect 4458 39136 4522 39140
rect 4538 39196 4602 39200
rect 4538 39140 4542 39196
rect 4542 39140 4598 39196
rect 4598 39140 4602 39196
rect 4538 39136 4602 39140
rect 4618 39196 4682 39200
rect 4618 39140 4622 39196
rect 4622 39140 4678 39196
rect 4678 39140 4682 39196
rect 4618 39136 4682 39140
rect 7805 39196 7869 39200
rect 7805 39140 7809 39196
rect 7809 39140 7865 39196
rect 7865 39140 7869 39196
rect 7805 39136 7869 39140
rect 7885 39196 7949 39200
rect 7885 39140 7889 39196
rect 7889 39140 7945 39196
rect 7945 39140 7949 39196
rect 7885 39136 7949 39140
rect 7965 39196 8029 39200
rect 7965 39140 7969 39196
rect 7969 39140 8025 39196
rect 8025 39140 8029 39196
rect 7965 39136 8029 39140
rect 8045 39196 8109 39200
rect 8045 39140 8049 39196
rect 8049 39140 8105 39196
rect 8105 39140 8109 39196
rect 8045 39136 8109 39140
rect 11232 39196 11296 39200
rect 11232 39140 11236 39196
rect 11236 39140 11292 39196
rect 11292 39140 11296 39196
rect 11232 39136 11296 39140
rect 11312 39196 11376 39200
rect 11312 39140 11316 39196
rect 11316 39140 11372 39196
rect 11372 39140 11376 39196
rect 11312 39136 11376 39140
rect 11392 39196 11456 39200
rect 11392 39140 11396 39196
rect 11396 39140 11452 39196
rect 11452 39140 11456 39196
rect 11392 39136 11456 39140
rect 11472 39196 11536 39200
rect 11472 39140 11476 39196
rect 11476 39140 11532 39196
rect 11532 39140 11536 39196
rect 11472 39136 11536 39140
rect 14659 39196 14723 39200
rect 14659 39140 14663 39196
rect 14663 39140 14719 39196
rect 14719 39140 14723 39196
rect 14659 39136 14723 39140
rect 14739 39196 14803 39200
rect 14739 39140 14743 39196
rect 14743 39140 14799 39196
rect 14799 39140 14803 39196
rect 14739 39136 14803 39140
rect 14819 39196 14883 39200
rect 14819 39140 14823 39196
rect 14823 39140 14879 39196
rect 14879 39140 14883 39196
rect 14819 39136 14883 39140
rect 14899 39196 14963 39200
rect 14899 39140 14903 39196
rect 14903 39140 14959 39196
rect 14959 39140 14963 39196
rect 14899 39136 14963 39140
rect 2665 38652 2729 38656
rect 2665 38596 2669 38652
rect 2669 38596 2725 38652
rect 2725 38596 2729 38652
rect 2665 38592 2729 38596
rect 2745 38652 2809 38656
rect 2745 38596 2749 38652
rect 2749 38596 2805 38652
rect 2805 38596 2809 38652
rect 2745 38592 2809 38596
rect 2825 38652 2889 38656
rect 2825 38596 2829 38652
rect 2829 38596 2885 38652
rect 2885 38596 2889 38652
rect 2825 38592 2889 38596
rect 2905 38652 2969 38656
rect 2905 38596 2909 38652
rect 2909 38596 2965 38652
rect 2965 38596 2969 38652
rect 2905 38592 2969 38596
rect 6092 38652 6156 38656
rect 6092 38596 6096 38652
rect 6096 38596 6152 38652
rect 6152 38596 6156 38652
rect 6092 38592 6156 38596
rect 6172 38652 6236 38656
rect 6172 38596 6176 38652
rect 6176 38596 6232 38652
rect 6232 38596 6236 38652
rect 6172 38592 6236 38596
rect 6252 38652 6316 38656
rect 6252 38596 6256 38652
rect 6256 38596 6312 38652
rect 6312 38596 6316 38652
rect 6252 38592 6316 38596
rect 6332 38652 6396 38656
rect 6332 38596 6336 38652
rect 6336 38596 6392 38652
rect 6392 38596 6396 38652
rect 6332 38592 6396 38596
rect 9519 38652 9583 38656
rect 9519 38596 9523 38652
rect 9523 38596 9579 38652
rect 9579 38596 9583 38652
rect 9519 38592 9583 38596
rect 9599 38652 9663 38656
rect 9599 38596 9603 38652
rect 9603 38596 9659 38652
rect 9659 38596 9663 38652
rect 9599 38592 9663 38596
rect 9679 38652 9743 38656
rect 9679 38596 9683 38652
rect 9683 38596 9739 38652
rect 9739 38596 9743 38652
rect 9679 38592 9743 38596
rect 9759 38652 9823 38656
rect 9759 38596 9763 38652
rect 9763 38596 9819 38652
rect 9819 38596 9823 38652
rect 9759 38592 9823 38596
rect 12946 38652 13010 38656
rect 12946 38596 12950 38652
rect 12950 38596 13006 38652
rect 13006 38596 13010 38652
rect 12946 38592 13010 38596
rect 13026 38652 13090 38656
rect 13026 38596 13030 38652
rect 13030 38596 13086 38652
rect 13086 38596 13090 38652
rect 13026 38592 13090 38596
rect 13106 38652 13170 38656
rect 13106 38596 13110 38652
rect 13110 38596 13166 38652
rect 13166 38596 13170 38652
rect 13106 38592 13170 38596
rect 13186 38652 13250 38656
rect 13186 38596 13190 38652
rect 13190 38596 13246 38652
rect 13246 38596 13250 38652
rect 13186 38592 13250 38596
rect 4378 38108 4442 38112
rect 4378 38052 4382 38108
rect 4382 38052 4438 38108
rect 4438 38052 4442 38108
rect 4378 38048 4442 38052
rect 4458 38108 4522 38112
rect 4458 38052 4462 38108
rect 4462 38052 4518 38108
rect 4518 38052 4522 38108
rect 4458 38048 4522 38052
rect 4538 38108 4602 38112
rect 4538 38052 4542 38108
rect 4542 38052 4598 38108
rect 4598 38052 4602 38108
rect 4538 38048 4602 38052
rect 4618 38108 4682 38112
rect 4618 38052 4622 38108
rect 4622 38052 4678 38108
rect 4678 38052 4682 38108
rect 4618 38048 4682 38052
rect 7805 38108 7869 38112
rect 7805 38052 7809 38108
rect 7809 38052 7865 38108
rect 7865 38052 7869 38108
rect 7805 38048 7869 38052
rect 7885 38108 7949 38112
rect 7885 38052 7889 38108
rect 7889 38052 7945 38108
rect 7945 38052 7949 38108
rect 7885 38048 7949 38052
rect 7965 38108 8029 38112
rect 7965 38052 7969 38108
rect 7969 38052 8025 38108
rect 8025 38052 8029 38108
rect 7965 38048 8029 38052
rect 8045 38108 8109 38112
rect 8045 38052 8049 38108
rect 8049 38052 8105 38108
rect 8105 38052 8109 38108
rect 8045 38048 8109 38052
rect 11232 38108 11296 38112
rect 11232 38052 11236 38108
rect 11236 38052 11292 38108
rect 11292 38052 11296 38108
rect 11232 38048 11296 38052
rect 11312 38108 11376 38112
rect 11312 38052 11316 38108
rect 11316 38052 11372 38108
rect 11372 38052 11376 38108
rect 11312 38048 11376 38052
rect 11392 38108 11456 38112
rect 11392 38052 11396 38108
rect 11396 38052 11452 38108
rect 11452 38052 11456 38108
rect 11392 38048 11456 38052
rect 11472 38108 11536 38112
rect 11472 38052 11476 38108
rect 11476 38052 11532 38108
rect 11532 38052 11536 38108
rect 11472 38048 11536 38052
rect 14659 38108 14723 38112
rect 14659 38052 14663 38108
rect 14663 38052 14719 38108
rect 14719 38052 14723 38108
rect 14659 38048 14723 38052
rect 14739 38108 14803 38112
rect 14739 38052 14743 38108
rect 14743 38052 14799 38108
rect 14799 38052 14803 38108
rect 14739 38048 14803 38052
rect 14819 38108 14883 38112
rect 14819 38052 14823 38108
rect 14823 38052 14879 38108
rect 14879 38052 14883 38108
rect 14819 38048 14883 38052
rect 14899 38108 14963 38112
rect 14899 38052 14903 38108
rect 14903 38052 14959 38108
rect 14959 38052 14963 38108
rect 14899 38048 14963 38052
rect 2665 37564 2729 37568
rect 2665 37508 2669 37564
rect 2669 37508 2725 37564
rect 2725 37508 2729 37564
rect 2665 37504 2729 37508
rect 2745 37564 2809 37568
rect 2745 37508 2749 37564
rect 2749 37508 2805 37564
rect 2805 37508 2809 37564
rect 2745 37504 2809 37508
rect 2825 37564 2889 37568
rect 2825 37508 2829 37564
rect 2829 37508 2885 37564
rect 2885 37508 2889 37564
rect 2825 37504 2889 37508
rect 2905 37564 2969 37568
rect 2905 37508 2909 37564
rect 2909 37508 2965 37564
rect 2965 37508 2969 37564
rect 2905 37504 2969 37508
rect 6092 37564 6156 37568
rect 6092 37508 6096 37564
rect 6096 37508 6152 37564
rect 6152 37508 6156 37564
rect 6092 37504 6156 37508
rect 6172 37564 6236 37568
rect 6172 37508 6176 37564
rect 6176 37508 6232 37564
rect 6232 37508 6236 37564
rect 6172 37504 6236 37508
rect 6252 37564 6316 37568
rect 6252 37508 6256 37564
rect 6256 37508 6312 37564
rect 6312 37508 6316 37564
rect 6252 37504 6316 37508
rect 6332 37564 6396 37568
rect 6332 37508 6336 37564
rect 6336 37508 6392 37564
rect 6392 37508 6396 37564
rect 6332 37504 6396 37508
rect 9519 37564 9583 37568
rect 9519 37508 9523 37564
rect 9523 37508 9579 37564
rect 9579 37508 9583 37564
rect 9519 37504 9583 37508
rect 9599 37564 9663 37568
rect 9599 37508 9603 37564
rect 9603 37508 9659 37564
rect 9659 37508 9663 37564
rect 9599 37504 9663 37508
rect 9679 37564 9743 37568
rect 9679 37508 9683 37564
rect 9683 37508 9739 37564
rect 9739 37508 9743 37564
rect 9679 37504 9743 37508
rect 9759 37564 9823 37568
rect 9759 37508 9763 37564
rect 9763 37508 9819 37564
rect 9819 37508 9823 37564
rect 9759 37504 9823 37508
rect 12946 37564 13010 37568
rect 12946 37508 12950 37564
rect 12950 37508 13006 37564
rect 13006 37508 13010 37564
rect 12946 37504 13010 37508
rect 13026 37564 13090 37568
rect 13026 37508 13030 37564
rect 13030 37508 13086 37564
rect 13086 37508 13090 37564
rect 13026 37504 13090 37508
rect 13106 37564 13170 37568
rect 13106 37508 13110 37564
rect 13110 37508 13166 37564
rect 13166 37508 13170 37564
rect 13106 37504 13170 37508
rect 13186 37564 13250 37568
rect 13186 37508 13190 37564
rect 13190 37508 13246 37564
rect 13246 37508 13250 37564
rect 13186 37504 13250 37508
rect 4378 37020 4442 37024
rect 4378 36964 4382 37020
rect 4382 36964 4438 37020
rect 4438 36964 4442 37020
rect 4378 36960 4442 36964
rect 4458 37020 4522 37024
rect 4458 36964 4462 37020
rect 4462 36964 4518 37020
rect 4518 36964 4522 37020
rect 4458 36960 4522 36964
rect 4538 37020 4602 37024
rect 4538 36964 4542 37020
rect 4542 36964 4598 37020
rect 4598 36964 4602 37020
rect 4538 36960 4602 36964
rect 4618 37020 4682 37024
rect 4618 36964 4622 37020
rect 4622 36964 4678 37020
rect 4678 36964 4682 37020
rect 4618 36960 4682 36964
rect 7805 37020 7869 37024
rect 7805 36964 7809 37020
rect 7809 36964 7865 37020
rect 7865 36964 7869 37020
rect 7805 36960 7869 36964
rect 7885 37020 7949 37024
rect 7885 36964 7889 37020
rect 7889 36964 7945 37020
rect 7945 36964 7949 37020
rect 7885 36960 7949 36964
rect 7965 37020 8029 37024
rect 7965 36964 7969 37020
rect 7969 36964 8025 37020
rect 8025 36964 8029 37020
rect 7965 36960 8029 36964
rect 8045 37020 8109 37024
rect 8045 36964 8049 37020
rect 8049 36964 8105 37020
rect 8105 36964 8109 37020
rect 8045 36960 8109 36964
rect 11232 37020 11296 37024
rect 11232 36964 11236 37020
rect 11236 36964 11292 37020
rect 11292 36964 11296 37020
rect 11232 36960 11296 36964
rect 11312 37020 11376 37024
rect 11312 36964 11316 37020
rect 11316 36964 11372 37020
rect 11372 36964 11376 37020
rect 11312 36960 11376 36964
rect 11392 37020 11456 37024
rect 11392 36964 11396 37020
rect 11396 36964 11452 37020
rect 11452 36964 11456 37020
rect 11392 36960 11456 36964
rect 11472 37020 11536 37024
rect 11472 36964 11476 37020
rect 11476 36964 11532 37020
rect 11532 36964 11536 37020
rect 11472 36960 11536 36964
rect 14659 37020 14723 37024
rect 14659 36964 14663 37020
rect 14663 36964 14719 37020
rect 14719 36964 14723 37020
rect 14659 36960 14723 36964
rect 14739 37020 14803 37024
rect 14739 36964 14743 37020
rect 14743 36964 14799 37020
rect 14799 36964 14803 37020
rect 14739 36960 14803 36964
rect 14819 37020 14883 37024
rect 14819 36964 14823 37020
rect 14823 36964 14879 37020
rect 14879 36964 14883 37020
rect 14819 36960 14883 36964
rect 14899 37020 14963 37024
rect 14899 36964 14903 37020
rect 14903 36964 14959 37020
rect 14959 36964 14963 37020
rect 14899 36960 14963 36964
rect 2665 36476 2729 36480
rect 2665 36420 2669 36476
rect 2669 36420 2725 36476
rect 2725 36420 2729 36476
rect 2665 36416 2729 36420
rect 2745 36476 2809 36480
rect 2745 36420 2749 36476
rect 2749 36420 2805 36476
rect 2805 36420 2809 36476
rect 2745 36416 2809 36420
rect 2825 36476 2889 36480
rect 2825 36420 2829 36476
rect 2829 36420 2885 36476
rect 2885 36420 2889 36476
rect 2825 36416 2889 36420
rect 2905 36476 2969 36480
rect 2905 36420 2909 36476
rect 2909 36420 2965 36476
rect 2965 36420 2969 36476
rect 2905 36416 2969 36420
rect 6092 36476 6156 36480
rect 6092 36420 6096 36476
rect 6096 36420 6152 36476
rect 6152 36420 6156 36476
rect 6092 36416 6156 36420
rect 6172 36476 6236 36480
rect 6172 36420 6176 36476
rect 6176 36420 6232 36476
rect 6232 36420 6236 36476
rect 6172 36416 6236 36420
rect 6252 36476 6316 36480
rect 6252 36420 6256 36476
rect 6256 36420 6312 36476
rect 6312 36420 6316 36476
rect 6252 36416 6316 36420
rect 6332 36476 6396 36480
rect 6332 36420 6336 36476
rect 6336 36420 6392 36476
rect 6392 36420 6396 36476
rect 6332 36416 6396 36420
rect 9519 36476 9583 36480
rect 9519 36420 9523 36476
rect 9523 36420 9579 36476
rect 9579 36420 9583 36476
rect 9519 36416 9583 36420
rect 9599 36476 9663 36480
rect 9599 36420 9603 36476
rect 9603 36420 9659 36476
rect 9659 36420 9663 36476
rect 9599 36416 9663 36420
rect 9679 36476 9743 36480
rect 9679 36420 9683 36476
rect 9683 36420 9739 36476
rect 9739 36420 9743 36476
rect 9679 36416 9743 36420
rect 9759 36476 9823 36480
rect 9759 36420 9763 36476
rect 9763 36420 9819 36476
rect 9819 36420 9823 36476
rect 9759 36416 9823 36420
rect 12946 36476 13010 36480
rect 12946 36420 12950 36476
rect 12950 36420 13006 36476
rect 13006 36420 13010 36476
rect 12946 36416 13010 36420
rect 13026 36476 13090 36480
rect 13026 36420 13030 36476
rect 13030 36420 13086 36476
rect 13086 36420 13090 36476
rect 13026 36416 13090 36420
rect 13106 36476 13170 36480
rect 13106 36420 13110 36476
rect 13110 36420 13166 36476
rect 13166 36420 13170 36476
rect 13106 36416 13170 36420
rect 13186 36476 13250 36480
rect 13186 36420 13190 36476
rect 13190 36420 13246 36476
rect 13246 36420 13250 36476
rect 13186 36416 13250 36420
rect 10548 36000 10612 36004
rect 10548 35944 10562 36000
rect 10562 35944 10612 36000
rect 10548 35940 10612 35944
rect 4378 35932 4442 35936
rect 4378 35876 4382 35932
rect 4382 35876 4438 35932
rect 4438 35876 4442 35932
rect 4378 35872 4442 35876
rect 4458 35932 4522 35936
rect 4458 35876 4462 35932
rect 4462 35876 4518 35932
rect 4518 35876 4522 35932
rect 4458 35872 4522 35876
rect 4538 35932 4602 35936
rect 4538 35876 4542 35932
rect 4542 35876 4598 35932
rect 4598 35876 4602 35932
rect 4538 35872 4602 35876
rect 4618 35932 4682 35936
rect 4618 35876 4622 35932
rect 4622 35876 4678 35932
rect 4678 35876 4682 35932
rect 4618 35872 4682 35876
rect 7805 35932 7869 35936
rect 7805 35876 7809 35932
rect 7809 35876 7865 35932
rect 7865 35876 7869 35932
rect 7805 35872 7869 35876
rect 7885 35932 7949 35936
rect 7885 35876 7889 35932
rect 7889 35876 7945 35932
rect 7945 35876 7949 35932
rect 7885 35872 7949 35876
rect 7965 35932 8029 35936
rect 7965 35876 7969 35932
rect 7969 35876 8025 35932
rect 8025 35876 8029 35932
rect 7965 35872 8029 35876
rect 8045 35932 8109 35936
rect 8045 35876 8049 35932
rect 8049 35876 8105 35932
rect 8105 35876 8109 35932
rect 8045 35872 8109 35876
rect 11232 35932 11296 35936
rect 11232 35876 11236 35932
rect 11236 35876 11292 35932
rect 11292 35876 11296 35932
rect 11232 35872 11296 35876
rect 11312 35932 11376 35936
rect 11312 35876 11316 35932
rect 11316 35876 11372 35932
rect 11372 35876 11376 35932
rect 11312 35872 11376 35876
rect 11392 35932 11456 35936
rect 11392 35876 11396 35932
rect 11396 35876 11452 35932
rect 11452 35876 11456 35932
rect 11392 35872 11456 35876
rect 11472 35932 11536 35936
rect 11472 35876 11476 35932
rect 11476 35876 11532 35932
rect 11532 35876 11536 35932
rect 11472 35872 11536 35876
rect 14659 35932 14723 35936
rect 14659 35876 14663 35932
rect 14663 35876 14719 35932
rect 14719 35876 14723 35932
rect 14659 35872 14723 35876
rect 14739 35932 14803 35936
rect 14739 35876 14743 35932
rect 14743 35876 14799 35932
rect 14799 35876 14803 35932
rect 14739 35872 14803 35876
rect 14819 35932 14883 35936
rect 14819 35876 14823 35932
rect 14823 35876 14879 35932
rect 14879 35876 14883 35932
rect 14819 35872 14883 35876
rect 14899 35932 14963 35936
rect 14899 35876 14903 35932
rect 14903 35876 14959 35932
rect 14959 35876 14963 35932
rect 14899 35872 14963 35876
rect 2665 35388 2729 35392
rect 2665 35332 2669 35388
rect 2669 35332 2725 35388
rect 2725 35332 2729 35388
rect 2665 35328 2729 35332
rect 2745 35388 2809 35392
rect 2745 35332 2749 35388
rect 2749 35332 2805 35388
rect 2805 35332 2809 35388
rect 2745 35328 2809 35332
rect 2825 35388 2889 35392
rect 2825 35332 2829 35388
rect 2829 35332 2885 35388
rect 2885 35332 2889 35388
rect 2825 35328 2889 35332
rect 2905 35388 2969 35392
rect 2905 35332 2909 35388
rect 2909 35332 2965 35388
rect 2965 35332 2969 35388
rect 2905 35328 2969 35332
rect 6092 35388 6156 35392
rect 6092 35332 6096 35388
rect 6096 35332 6152 35388
rect 6152 35332 6156 35388
rect 6092 35328 6156 35332
rect 6172 35388 6236 35392
rect 6172 35332 6176 35388
rect 6176 35332 6232 35388
rect 6232 35332 6236 35388
rect 6172 35328 6236 35332
rect 6252 35388 6316 35392
rect 6252 35332 6256 35388
rect 6256 35332 6312 35388
rect 6312 35332 6316 35388
rect 6252 35328 6316 35332
rect 6332 35388 6396 35392
rect 6332 35332 6336 35388
rect 6336 35332 6392 35388
rect 6392 35332 6396 35388
rect 6332 35328 6396 35332
rect 9519 35388 9583 35392
rect 9519 35332 9523 35388
rect 9523 35332 9579 35388
rect 9579 35332 9583 35388
rect 9519 35328 9583 35332
rect 9599 35388 9663 35392
rect 9599 35332 9603 35388
rect 9603 35332 9659 35388
rect 9659 35332 9663 35388
rect 9599 35328 9663 35332
rect 9679 35388 9743 35392
rect 9679 35332 9683 35388
rect 9683 35332 9739 35388
rect 9739 35332 9743 35388
rect 9679 35328 9743 35332
rect 9759 35388 9823 35392
rect 9759 35332 9763 35388
rect 9763 35332 9819 35388
rect 9819 35332 9823 35388
rect 9759 35328 9823 35332
rect 12946 35388 13010 35392
rect 12946 35332 12950 35388
rect 12950 35332 13006 35388
rect 13006 35332 13010 35388
rect 12946 35328 13010 35332
rect 13026 35388 13090 35392
rect 13026 35332 13030 35388
rect 13030 35332 13086 35388
rect 13086 35332 13090 35388
rect 13026 35328 13090 35332
rect 13106 35388 13170 35392
rect 13106 35332 13110 35388
rect 13110 35332 13166 35388
rect 13166 35332 13170 35388
rect 13106 35328 13170 35332
rect 13186 35388 13250 35392
rect 13186 35332 13190 35388
rect 13190 35332 13246 35388
rect 13246 35332 13250 35388
rect 13186 35328 13250 35332
rect 4378 34844 4442 34848
rect 4378 34788 4382 34844
rect 4382 34788 4438 34844
rect 4438 34788 4442 34844
rect 4378 34784 4442 34788
rect 4458 34844 4522 34848
rect 4458 34788 4462 34844
rect 4462 34788 4518 34844
rect 4518 34788 4522 34844
rect 4458 34784 4522 34788
rect 4538 34844 4602 34848
rect 4538 34788 4542 34844
rect 4542 34788 4598 34844
rect 4598 34788 4602 34844
rect 4538 34784 4602 34788
rect 4618 34844 4682 34848
rect 4618 34788 4622 34844
rect 4622 34788 4678 34844
rect 4678 34788 4682 34844
rect 4618 34784 4682 34788
rect 7805 34844 7869 34848
rect 7805 34788 7809 34844
rect 7809 34788 7865 34844
rect 7865 34788 7869 34844
rect 7805 34784 7869 34788
rect 7885 34844 7949 34848
rect 7885 34788 7889 34844
rect 7889 34788 7945 34844
rect 7945 34788 7949 34844
rect 7885 34784 7949 34788
rect 7965 34844 8029 34848
rect 7965 34788 7969 34844
rect 7969 34788 8025 34844
rect 8025 34788 8029 34844
rect 7965 34784 8029 34788
rect 8045 34844 8109 34848
rect 8045 34788 8049 34844
rect 8049 34788 8105 34844
rect 8105 34788 8109 34844
rect 8045 34784 8109 34788
rect 11232 34844 11296 34848
rect 11232 34788 11236 34844
rect 11236 34788 11292 34844
rect 11292 34788 11296 34844
rect 11232 34784 11296 34788
rect 11312 34844 11376 34848
rect 11312 34788 11316 34844
rect 11316 34788 11372 34844
rect 11372 34788 11376 34844
rect 11312 34784 11376 34788
rect 11392 34844 11456 34848
rect 11392 34788 11396 34844
rect 11396 34788 11452 34844
rect 11452 34788 11456 34844
rect 11392 34784 11456 34788
rect 11472 34844 11536 34848
rect 11472 34788 11476 34844
rect 11476 34788 11532 34844
rect 11532 34788 11536 34844
rect 11472 34784 11536 34788
rect 14659 34844 14723 34848
rect 14659 34788 14663 34844
rect 14663 34788 14719 34844
rect 14719 34788 14723 34844
rect 14659 34784 14723 34788
rect 14739 34844 14803 34848
rect 14739 34788 14743 34844
rect 14743 34788 14799 34844
rect 14799 34788 14803 34844
rect 14739 34784 14803 34788
rect 14819 34844 14883 34848
rect 14819 34788 14823 34844
rect 14823 34788 14879 34844
rect 14879 34788 14883 34844
rect 14819 34784 14883 34788
rect 14899 34844 14963 34848
rect 14899 34788 14903 34844
rect 14903 34788 14959 34844
rect 14959 34788 14963 34844
rect 14899 34784 14963 34788
rect 2665 34300 2729 34304
rect 2665 34244 2669 34300
rect 2669 34244 2725 34300
rect 2725 34244 2729 34300
rect 2665 34240 2729 34244
rect 2745 34300 2809 34304
rect 2745 34244 2749 34300
rect 2749 34244 2805 34300
rect 2805 34244 2809 34300
rect 2745 34240 2809 34244
rect 2825 34300 2889 34304
rect 2825 34244 2829 34300
rect 2829 34244 2885 34300
rect 2885 34244 2889 34300
rect 2825 34240 2889 34244
rect 2905 34300 2969 34304
rect 2905 34244 2909 34300
rect 2909 34244 2965 34300
rect 2965 34244 2969 34300
rect 2905 34240 2969 34244
rect 6092 34300 6156 34304
rect 6092 34244 6096 34300
rect 6096 34244 6152 34300
rect 6152 34244 6156 34300
rect 6092 34240 6156 34244
rect 6172 34300 6236 34304
rect 6172 34244 6176 34300
rect 6176 34244 6232 34300
rect 6232 34244 6236 34300
rect 6172 34240 6236 34244
rect 6252 34300 6316 34304
rect 6252 34244 6256 34300
rect 6256 34244 6312 34300
rect 6312 34244 6316 34300
rect 6252 34240 6316 34244
rect 6332 34300 6396 34304
rect 6332 34244 6336 34300
rect 6336 34244 6392 34300
rect 6392 34244 6396 34300
rect 6332 34240 6396 34244
rect 9519 34300 9583 34304
rect 9519 34244 9523 34300
rect 9523 34244 9579 34300
rect 9579 34244 9583 34300
rect 9519 34240 9583 34244
rect 9599 34300 9663 34304
rect 9599 34244 9603 34300
rect 9603 34244 9659 34300
rect 9659 34244 9663 34300
rect 9599 34240 9663 34244
rect 9679 34300 9743 34304
rect 9679 34244 9683 34300
rect 9683 34244 9739 34300
rect 9739 34244 9743 34300
rect 9679 34240 9743 34244
rect 9759 34300 9823 34304
rect 9759 34244 9763 34300
rect 9763 34244 9819 34300
rect 9819 34244 9823 34300
rect 9759 34240 9823 34244
rect 12946 34300 13010 34304
rect 12946 34244 12950 34300
rect 12950 34244 13006 34300
rect 13006 34244 13010 34300
rect 12946 34240 13010 34244
rect 13026 34300 13090 34304
rect 13026 34244 13030 34300
rect 13030 34244 13086 34300
rect 13086 34244 13090 34300
rect 13026 34240 13090 34244
rect 13106 34300 13170 34304
rect 13106 34244 13110 34300
rect 13110 34244 13166 34300
rect 13166 34244 13170 34300
rect 13106 34240 13170 34244
rect 13186 34300 13250 34304
rect 13186 34244 13190 34300
rect 13190 34244 13246 34300
rect 13246 34244 13250 34300
rect 13186 34240 13250 34244
rect 11652 33900 11716 33964
rect 4378 33756 4442 33760
rect 4378 33700 4382 33756
rect 4382 33700 4438 33756
rect 4438 33700 4442 33756
rect 4378 33696 4442 33700
rect 4458 33756 4522 33760
rect 4458 33700 4462 33756
rect 4462 33700 4518 33756
rect 4518 33700 4522 33756
rect 4458 33696 4522 33700
rect 4538 33756 4602 33760
rect 4538 33700 4542 33756
rect 4542 33700 4598 33756
rect 4598 33700 4602 33756
rect 4538 33696 4602 33700
rect 4618 33756 4682 33760
rect 4618 33700 4622 33756
rect 4622 33700 4678 33756
rect 4678 33700 4682 33756
rect 4618 33696 4682 33700
rect 7805 33756 7869 33760
rect 7805 33700 7809 33756
rect 7809 33700 7865 33756
rect 7865 33700 7869 33756
rect 7805 33696 7869 33700
rect 7885 33756 7949 33760
rect 7885 33700 7889 33756
rect 7889 33700 7945 33756
rect 7945 33700 7949 33756
rect 7885 33696 7949 33700
rect 7965 33756 8029 33760
rect 7965 33700 7969 33756
rect 7969 33700 8025 33756
rect 8025 33700 8029 33756
rect 7965 33696 8029 33700
rect 8045 33756 8109 33760
rect 8045 33700 8049 33756
rect 8049 33700 8105 33756
rect 8105 33700 8109 33756
rect 8045 33696 8109 33700
rect 11232 33756 11296 33760
rect 11232 33700 11236 33756
rect 11236 33700 11292 33756
rect 11292 33700 11296 33756
rect 11232 33696 11296 33700
rect 11312 33756 11376 33760
rect 11312 33700 11316 33756
rect 11316 33700 11372 33756
rect 11372 33700 11376 33756
rect 11312 33696 11376 33700
rect 11392 33756 11456 33760
rect 11392 33700 11396 33756
rect 11396 33700 11452 33756
rect 11452 33700 11456 33756
rect 11392 33696 11456 33700
rect 11472 33756 11536 33760
rect 11472 33700 11476 33756
rect 11476 33700 11532 33756
rect 11532 33700 11536 33756
rect 11472 33696 11536 33700
rect 14659 33756 14723 33760
rect 14659 33700 14663 33756
rect 14663 33700 14719 33756
rect 14719 33700 14723 33756
rect 14659 33696 14723 33700
rect 14739 33756 14803 33760
rect 14739 33700 14743 33756
rect 14743 33700 14799 33756
rect 14799 33700 14803 33756
rect 14739 33696 14803 33700
rect 14819 33756 14883 33760
rect 14819 33700 14823 33756
rect 14823 33700 14879 33756
rect 14879 33700 14883 33756
rect 14819 33696 14883 33700
rect 14899 33756 14963 33760
rect 14899 33700 14903 33756
rect 14903 33700 14959 33756
rect 14959 33700 14963 33756
rect 14899 33696 14963 33700
rect 13492 33628 13556 33692
rect 8892 33220 8956 33284
rect 2665 33212 2729 33216
rect 2665 33156 2669 33212
rect 2669 33156 2725 33212
rect 2725 33156 2729 33212
rect 2665 33152 2729 33156
rect 2745 33212 2809 33216
rect 2745 33156 2749 33212
rect 2749 33156 2805 33212
rect 2805 33156 2809 33212
rect 2745 33152 2809 33156
rect 2825 33212 2889 33216
rect 2825 33156 2829 33212
rect 2829 33156 2885 33212
rect 2885 33156 2889 33212
rect 2825 33152 2889 33156
rect 2905 33212 2969 33216
rect 2905 33156 2909 33212
rect 2909 33156 2965 33212
rect 2965 33156 2969 33212
rect 2905 33152 2969 33156
rect 6092 33212 6156 33216
rect 6092 33156 6096 33212
rect 6096 33156 6152 33212
rect 6152 33156 6156 33212
rect 6092 33152 6156 33156
rect 6172 33212 6236 33216
rect 6172 33156 6176 33212
rect 6176 33156 6232 33212
rect 6232 33156 6236 33212
rect 6172 33152 6236 33156
rect 6252 33212 6316 33216
rect 6252 33156 6256 33212
rect 6256 33156 6312 33212
rect 6312 33156 6316 33212
rect 6252 33152 6316 33156
rect 6332 33212 6396 33216
rect 6332 33156 6336 33212
rect 6336 33156 6392 33212
rect 6392 33156 6396 33212
rect 6332 33152 6396 33156
rect 9519 33212 9583 33216
rect 9519 33156 9523 33212
rect 9523 33156 9579 33212
rect 9579 33156 9583 33212
rect 9519 33152 9583 33156
rect 9599 33212 9663 33216
rect 9599 33156 9603 33212
rect 9603 33156 9659 33212
rect 9659 33156 9663 33212
rect 9599 33152 9663 33156
rect 9679 33212 9743 33216
rect 9679 33156 9683 33212
rect 9683 33156 9739 33212
rect 9739 33156 9743 33212
rect 9679 33152 9743 33156
rect 9759 33212 9823 33216
rect 9759 33156 9763 33212
rect 9763 33156 9819 33212
rect 9819 33156 9823 33212
rect 9759 33152 9823 33156
rect 12946 33212 13010 33216
rect 12946 33156 12950 33212
rect 12950 33156 13006 33212
rect 13006 33156 13010 33212
rect 12946 33152 13010 33156
rect 13026 33212 13090 33216
rect 13026 33156 13030 33212
rect 13030 33156 13086 33212
rect 13086 33156 13090 33212
rect 13026 33152 13090 33156
rect 13106 33212 13170 33216
rect 13106 33156 13110 33212
rect 13110 33156 13166 33212
rect 13166 33156 13170 33212
rect 13106 33152 13170 33156
rect 13186 33212 13250 33216
rect 13186 33156 13190 33212
rect 13190 33156 13246 33212
rect 13246 33156 13250 33212
rect 13186 33152 13250 33156
rect 12756 32676 12820 32740
rect 4378 32668 4442 32672
rect 4378 32612 4382 32668
rect 4382 32612 4438 32668
rect 4438 32612 4442 32668
rect 4378 32608 4442 32612
rect 4458 32668 4522 32672
rect 4458 32612 4462 32668
rect 4462 32612 4518 32668
rect 4518 32612 4522 32668
rect 4458 32608 4522 32612
rect 4538 32668 4602 32672
rect 4538 32612 4542 32668
rect 4542 32612 4598 32668
rect 4598 32612 4602 32668
rect 4538 32608 4602 32612
rect 4618 32668 4682 32672
rect 4618 32612 4622 32668
rect 4622 32612 4678 32668
rect 4678 32612 4682 32668
rect 4618 32608 4682 32612
rect 7805 32668 7869 32672
rect 7805 32612 7809 32668
rect 7809 32612 7865 32668
rect 7865 32612 7869 32668
rect 7805 32608 7869 32612
rect 7885 32668 7949 32672
rect 7885 32612 7889 32668
rect 7889 32612 7945 32668
rect 7945 32612 7949 32668
rect 7885 32608 7949 32612
rect 7965 32668 8029 32672
rect 7965 32612 7969 32668
rect 7969 32612 8025 32668
rect 8025 32612 8029 32668
rect 7965 32608 8029 32612
rect 8045 32668 8109 32672
rect 8045 32612 8049 32668
rect 8049 32612 8105 32668
rect 8105 32612 8109 32668
rect 8045 32608 8109 32612
rect 11232 32668 11296 32672
rect 11232 32612 11236 32668
rect 11236 32612 11292 32668
rect 11292 32612 11296 32668
rect 11232 32608 11296 32612
rect 11312 32668 11376 32672
rect 11312 32612 11316 32668
rect 11316 32612 11372 32668
rect 11372 32612 11376 32668
rect 11312 32608 11376 32612
rect 11392 32668 11456 32672
rect 11392 32612 11396 32668
rect 11396 32612 11452 32668
rect 11452 32612 11456 32668
rect 11392 32608 11456 32612
rect 11472 32668 11536 32672
rect 11472 32612 11476 32668
rect 11476 32612 11532 32668
rect 11532 32612 11536 32668
rect 11472 32608 11536 32612
rect 14659 32668 14723 32672
rect 14659 32612 14663 32668
rect 14663 32612 14719 32668
rect 14719 32612 14723 32668
rect 14659 32608 14723 32612
rect 14739 32668 14803 32672
rect 14739 32612 14743 32668
rect 14743 32612 14799 32668
rect 14799 32612 14803 32668
rect 14739 32608 14803 32612
rect 14819 32668 14883 32672
rect 14819 32612 14823 32668
rect 14823 32612 14879 32668
rect 14879 32612 14883 32668
rect 14819 32608 14883 32612
rect 14899 32668 14963 32672
rect 14899 32612 14903 32668
rect 14903 32612 14959 32668
rect 14959 32612 14963 32668
rect 14899 32608 14963 32612
rect 12572 32600 12636 32604
rect 12572 32544 12622 32600
rect 12622 32544 12636 32600
rect 12572 32540 12636 32544
rect 2665 32124 2729 32128
rect 2665 32068 2669 32124
rect 2669 32068 2725 32124
rect 2725 32068 2729 32124
rect 2665 32064 2729 32068
rect 2745 32124 2809 32128
rect 2745 32068 2749 32124
rect 2749 32068 2805 32124
rect 2805 32068 2809 32124
rect 2745 32064 2809 32068
rect 2825 32124 2889 32128
rect 2825 32068 2829 32124
rect 2829 32068 2885 32124
rect 2885 32068 2889 32124
rect 2825 32064 2889 32068
rect 2905 32124 2969 32128
rect 2905 32068 2909 32124
rect 2909 32068 2965 32124
rect 2965 32068 2969 32124
rect 2905 32064 2969 32068
rect 6092 32124 6156 32128
rect 6092 32068 6096 32124
rect 6096 32068 6152 32124
rect 6152 32068 6156 32124
rect 6092 32064 6156 32068
rect 6172 32124 6236 32128
rect 6172 32068 6176 32124
rect 6176 32068 6232 32124
rect 6232 32068 6236 32124
rect 6172 32064 6236 32068
rect 6252 32124 6316 32128
rect 6252 32068 6256 32124
rect 6256 32068 6312 32124
rect 6312 32068 6316 32124
rect 6252 32064 6316 32068
rect 6332 32124 6396 32128
rect 6332 32068 6336 32124
rect 6336 32068 6392 32124
rect 6392 32068 6396 32124
rect 6332 32064 6396 32068
rect 9519 32124 9583 32128
rect 9519 32068 9523 32124
rect 9523 32068 9579 32124
rect 9579 32068 9583 32124
rect 9519 32064 9583 32068
rect 9599 32124 9663 32128
rect 9599 32068 9603 32124
rect 9603 32068 9659 32124
rect 9659 32068 9663 32124
rect 9599 32064 9663 32068
rect 9679 32124 9743 32128
rect 9679 32068 9683 32124
rect 9683 32068 9739 32124
rect 9739 32068 9743 32124
rect 9679 32064 9743 32068
rect 9759 32124 9823 32128
rect 9759 32068 9763 32124
rect 9763 32068 9819 32124
rect 9819 32068 9823 32124
rect 9759 32064 9823 32068
rect 12946 32124 13010 32128
rect 12946 32068 12950 32124
rect 12950 32068 13006 32124
rect 13006 32068 13010 32124
rect 12946 32064 13010 32068
rect 13026 32124 13090 32128
rect 13026 32068 13030 32124
rect 13030 32068 13086 32124
rect 13086 32068 13090 32124
rect 13026 32064 13090 32068
rect 13106 32124 13170 32128
rect 13106 32068 13110 32124
rect 13110 32068 13166 32124
rect 13166 32068 13170 32124
rect 13106 32064 13170 32068
rect 13186 32124 13250 32128
rect 13186 32068 13190 32124
rect 13190 32068 13246 32124
rect 13246 32068 13250 32124
rect 13186 32064 13250 32068
rect 7236 31860 7300 31924
rect 14044 31724 14108 31788
rect 4378 31580 4442 31584
rect 4378 31524 4382 31580
rect 4382 31524 4438 31580
rect 4438 31524 4442 31580
rect 4378 31520 4442 31524
rect 4458 31580 4522 31584
rect 4458 31524 4462 31580
rect 4462 31524 4518 31580
rect 4518 31524 4522 31580
rect 4458 31520 4522 31524
rect 4538 31580 4602 31584
rect 4538 31524 4542 31580
rect 4542 31524 4598 31580
rect 4598 31524 4602 31580
rect 4538 31520 4602 31524
rect 4618 31580 4682 31584
rect 4618 31524 4622 31580
rect 4622 31524 4678 31580
rect 4678 31524 4682 31580
rect 4618 31520 4682 31524
rect 7805 31580 7869 31584
rect 7805 31524 7809 31580
rect 7809 31524 7865 31580
rect 7865 31524 7869 31580
rect 7805 31520 7869 31524
rect 7885 31580 7949 31584
rect 7885 31524 7889 31580
rect 7889 31524 7945 31580
rect 7945 31524 7949 31580
rect 7885 31520 7949 31524
rect 7965 31580 8029 31584
rect 7965 31524 7969 31580
rect 7969 31524 8025 31580
rect 8025 31524 8029 31580
rect 7965 31520 8029 31524
rect 8045 31580 8109 31584
rect 8045 31524 8049 31580
rect 8049 31524 8105 31580
rect 8105 31524 8109 31580
rect 8045 31520 8109 31524
rect 11232 31580 11296 31584
rect 11232 31524 11236 31580
rect 11236 31524 11292 31580
rect 11292 31524 11296 31580
rect 11232 31520 11296 31524
rect 11312 31580 11376 31584
rect 11312 31524 11316 31580
rect 11316 31524 11372 31580
rect 11372 31524 11376 31580
rect 11312 31520 11376 31524
rect 11392 31580 11456 31584
rect 11392 31524 11396 31580
rect 11396 31524 11452 31580
rect 11452 31524 11456 31580
rect 11392 31520 11456 31524
rect 11472 31580 11536 31584
rect 11472 31524 11476 31580
rect 11476 31524 11532 31580
rect 11532 31524 11536 31580
rect 11472 31520 11536 31524
rect 14659 31580 14723 31584
rect 14659 31524 14663 31580
rect 14663 31524 14719 31580
rect 14719 31524 14723 31580
rect 14659 31520 14723 31524
rect 14739 31580 14803 31584
rect 14739 31524 14743 31580
rect 14743 31524 14799 31580
rect 14799 31524 14803 31580
rect 14739 31520 14803 31524
rect 14819 31580 14883 31584
rect 14819 31524 14823 31580
rect 14823 31524 14879 31580
rect 14879 31524 14883 31580
rect 14819 31520 14883 31524
rect 14899 31580 14963 31584
rect 14899 31524 14903 31580
rect 14903 31524 14959 31580
rect 14959 31524 14963 31580
rect 14899 31520 14963 31524
rect 2665 31036 2729 31040
rect 2665 30980 2669 31036
rect 2669 30980 2725 31036
rect 2725 30980 2729 31036
rect 2665 30976 2729 30980
rect 2745 31036 2809 31040
rect 2745 30980 2749 31036
rect 2749 30980 2805 31036
rect 2805 30980 2809 31036
rect 2745 30976 2809 30980
rect 2825 31036 2889 31040
rect 2825 30980 2829 31036
rect 2829 30980 2885 31036
rect 2885 30980 2889 31036
rect 2825 30976 2889 30980
rect 2905 31036 2969 31040
rect 2905 30980 2909 31036
rect 2909 30980 2965 31036
rect 2965 30980 2969 31036
rect 2905 30976 2969 30980
rect 6092 31036 6156 31040
rect 6092 30980 6096 31036
rect 6096 30980 6152 31036
rect 6152 30980 6156 31036
rect 6092 30976 6156 30980
rect 6172 31036 6236 31040
rect 6172 30980 6176 31036
rect 6176 30980 6232 31036
rect 6232 30980 6236 31036
rect 6172 30976 6236 30980
rect 6252 31036 6316 31040
rect 6252 30980 6256 31036
rect 6256 30980 6312 31036
rect 6312 30980 6316 31036
rect 6252 30976 6316 30980
rect 6332 31036 6396 31040
rect 6332 30980 6336 31036
rect 6336 30980 6392 31036
rect 6392 30980 6396 31036
rect 6332 30976 6396 30980
rect 9519 31036 9583 31040
rect 9519 30980 9523 31036
rect 9523 30980 9579 31036
rect 9579 30980 9583 31036
rect 9519 30976 9583 30980
rect 9599 31036 9663 31040
rect 9599 30980 9603 31036
rect 9603 30980 9659 31036
rect 9659 30980 9663 31036
rect 9599 30976 9663 30980
rect 9679 31036 9743 31040
rect 9679 30980 9683 31036
rect 9683 30980 9739 31036
rect 9739 30980 9743 31036
rect 9679 30976 9743 30980
rect 9759 31036 9823 31040
rect 9759 30980 9763 31036
rect 9763 30980 9819 31036
rect 9819 30980 9823 31036
rect 9759 30976 9823 30980
rect 12946 31036 13010 31040
rect 12946 30980 12950 31036
rect 12950 30980 13006 31036
rect 13006 30980 13010 31036
rect 12946 30976 13010 30980
rect 13026 31036 13090 31040
rect 13026 30980 13030 31036
rect 13030 30980 13086 31036
rect 13086 30980 13090 31036
rect 13026 30976 13090 30980
rect 13106 31036 13170 31040
rect 13106 30980 13110 31036
rect 13110 30980 13166 31036
rect 13166 30980 13170 31036
rect 13106 30976 13170 30980
rect 13186 31036 13250 31040
rect 13186 30980 13190 31036
rect 13190 30980 13246 31036
rect 13246 30980 13250 31036
rect 13186 30976 13250 30980
rect 9076 30772 9140 30836
rect 10732 30636 10796 30700
rect 4378 30492 4442 30496
rect 4378 30436 4382 30492
rect 4382 30436 4438 30492
rect 4438 30436 4442 30492
rect 4378 30432 4442 30436
rect 4458 30492 4522 30496
rect 4458 30436 4462 30492
rect 4462 30436 4518 30492
rect 4518 30436 4522 30492
rect 4458 30432 4522 30436
rect 4538 30492 4602 30496
rect 4538 30436 4542 30492
rect 4542 30436 4598 30492
rect 4598 30436 4602 30492
rect 4538 30432 4602 30436
rect 4618 30492 4682 30496
rect 4618 30436 4622 30492
rect 4622 30436 4678 30492
rect 4678 30436 4682 30492
rect 4618 30432 4682 30436
rect 7805 30492 7869 30496
rect 7805 30436 7809 30492
rect 7809 30436 7865 30492
rect 7865 30436 7869 30492
rect 7805 30432 7869 30436
rect 7885 30492 7949 30496
rect 7885 30436 7889 30492
rect 7889 30436 7945 30492
rect 7945 30436 7949 30492
rect 7885 30432 7949 30436
rect 7965 30492 8029 30496
rect 7965 30436 7969 30492
rect 7969 30436 8025 30492
rect 8025 30436 8029 30492
rect 7965 30432 8029 30436
rect 8045 30492 8109 30496
rect 8045 30436 8049 30492
rect 8049 30436 8105 30492
rect 8105 30436 8109 30492
rect 8045 30432 8109 30436
rect 11232 30492 11296 30496
rect 11232 30436 11236 30492
rect 11236 30436 11292 30492
rect 11292 30436 11296 30492
rect 11232 30432 11296 30436
rect 11312 30492 11376 30496
rect 11312 30436 11316 30492
rect 11316 30436 11372 30492
rect 11372 30436 11376 30492
rect 11312 30432 11376 30436
rect 11392 30492 11456 30496
rect 11392 30436 11396 30492
rect 11396 30436 11452 30492
rect 11452 30436 11456 30492
rect 11392 30432 11456 30436
rect 11472 30492 11536 30496
rect 11472 30436 11476 30492
rect 11476 30436 11532 30492
rect 11532 30436 11536 30492
rect 11472 30432 11536 30436
rect 14659 30492 14723 30496
rect 14659 30436 14663 30492
rect 14663 30436 14719 30492
rect 14719 30436 14723 30492
rect 14659 30432 14723 30436
rect 14739 30492 14803 30496
rect 14739 30436 14743 30492
rect 14743 30436 14799 30492
rect 14799 30436 14803 30492
rect 14739 30432 14803 30436
rect 14819 30492 14883 30496
rect 14819 30436 14823 30492
rect 14823 30436 14879 30492
rect 14879 30436 14883 30492
rect 14819 30432 14883 30436
rect 14899 30492 14963 30496
rect 14899 30436 14903 30492
rect 14903 30436 14959 30492
rect 14959 30436 14963 30492
rect 14899 30432 14963 30436
rect 12572 30092 12636 30156
rect 2665 29948 2729 29952
rect 2665 29892 2669 29948
rect 2669 29892 2725 29948
rect 2725 29892 2729 29948
rect 2665 29888 2729 29892
rect 2745 29948 2809 29952
rect 2745 29892 2749 29948
rect 2749 29892 2805 29948
rect 2805 29892 2809 29948
rect 2745 29888 2809 29892
rect 2825 29948 2889 29952
rect 2825 29892 2829 29948
rect 2829 29892 2885 29948
rect 2885 29892 2889 29948
rect 2825 29888 2889 29892
rect 2905 29948 2969 29952
rect 2905 29892 2909 29948
rect 2909 29892 2965 29948
rect 2965 29892 2969 29948
rect 2905 29888 2969 29892
rect 6092 29948 6156 29952
rect 6092 29892 6096 29948
rect 6096 29892 6152 29948
rect 6152 29892 6156 29948
rect 6092 29888 6156 29892
rect 6172 29948 6236 29952
rect 6172 29892 6176 29948
rect 6176 29892 6232 29948
rect 6232 29892 6236 29948
rect 6172 29888 6236 29892
rect 6252 29948 6316 29952
rect 6252 29892 6256 29948
rect 6256 29892 6312 29948
rect 6312 29892 6316 29948
rect 6252 29888 6316 29892
rect 6332 29948 6396 29952
rect 6332 29892 6336 29948
rect 6336 29892 6392 29948
rect 6392 29892 6396 29948
rect 6332 29888 6396 29892
rect 9519 29948 9583 29952
rect 9519 29892 9523 29948
rect 9523 29892 9579 29948
rect 9579 29892 9583 29948
rect 9519 29888 9583 29892
rect 9599 29948 9663 29952
rect 9599 29892 9603 29948
rect 9603 29892 9659 29948
rect 9659 29892 9663 29948
rect 9599 29888 9663 29892
rect 9679 29948 9743 29952
rect 9679 29892 9683 29948
rect 9683 29892 9739 29948
rect 9739 29892 9743 29948
rect 9679 29888 9743 29892
rect 9759 29948 9823 29952
rect 9759 29892 9763 29948
rect 9763 29892 9819 29948
rect 9819 29892 9823 29948
rect 9759 29888 9823 29892
rect 12946 29948 13010 29952
rect 12946 29892 12950 29948
rect 12950 29892 13006 29948
rect 13006 29892 13010 29948
rect 12946 29888 13010 29892
rect 13026 29948 13090 29952
rect 13026 29892 13030 29948
rect 13030 29892 13086 29948
rect 13086 29892 13090 29948
rect 13026 29888 13090 29892
rect 13106 29948 13170 29952
rect 13106 29892 13110 29948
rect 13110 29892 13166 29948
rect 13166 29892 13170 29948
rect 13106 29888 13170 29892
rect 13186 29948 13250 29952
rect 13186 29892 13190 29948
rect 13190 29892 13246 29948
rect 13246 29892 13250 29948
rect 13186 29888 13250 29892
rect 12756 29820 12820 29884
rect 10732 29548 10796 29612
rect 4378 29404 4442 29408
rect 4378 29348 4382 29404
rect 4382 29348 4438 29404
rect 4438 29348 4442 29404
rect 4378 29344 4442 29348
rect 4458 29404 4522 29408
rect 4458 29348 4462 29404
rect 4462 29348 4518 29404
rect 4518 29348 4522 29404
rect 4458 29344 4522 29348
rect 4538 29404 4602 29408
rect 4538 29348 4542 29404
rect 4542 29348 4598 29404
rect 4598 29348 4602 29404
rect 4538 29344 4602 29348
rect 4618 29404 4682 29408
rect 4618 29348 4622 29404
rect 4622 29348 4678 29404
rect 4678 29348 4682 29404
rect 4618 29344 4682 29348
rect 7805 29404 7869 29408
rect 7805 29348 7809 29404
rect 7809 29348 7865 29404
rect 7865 29348 7869 29404
rect 7805 29344 7869 29348
rect 7885 29404 7949 29408
rect 7885 29348 7889 29404
rect 7889 29348 7945 29404
rect 7945 29348 7949 29404
rect 7885 29344 7949 29348
rect 7965 29404 8029 29408
rect 7965 29348 7969 29404
rect 7969 29348 8025 29404
rect 8025 29348 8029 29404
rect 7965 29344 8029 29348
rect 8045 29404 8109 29408
rect 8045 29348 8049 29404
rect 8049 29348 8105 29404
rect 8105 29348 8109 29404
rect 8045 29344 8109 29348
rect 11232 29404 11296 29408
rect 11232 29348 11236 29404
rect 11236 29348 11292 29404
rect 11292 29348 11296 29404
rect 11232 29344 11296 29348
rect 11312 29404 11376 29408
rect 11312 29348 11316 29404
rect 11316 29348 11372 29404
rect 11372 29348 11376 29404
rect 11312 29344 11376 29348
rect 11392 29404 11456 29408
rect 11392 29348 11396 29404
rect 11396 29348 11452 29404
rect 11452 29348 11456 29404
rect 11392 29344 11456 29348
rect 11472 29404 11536 29408
rect 11472 29348 11476 29404
rect 11476 29348 11532 29404
rect 11532 29348 11536 29404
rect 11472 29344 11536 29348
rect 14659 29404 14723 29408
rect 14659 29348 14663 29404
rect 14663 29348 14719 29404
rect 14719 29348 14723 29404
rect 14659 29344 14723 29348
rect 14739 29404 14803 29408
rect 14739 29348 14743 29404
rect 14743 29348 14799 29404
rect 14799 29348 14803 29404
rect 14739 29344 14803 29348
rect 14819 29404 14883 29408
rect 14819 29348 14823 29404
rect 14823 29348 14879 29404
rect 14879 29348 14883 29404
rect 14819 29344 14883 29348
rect 14899 29404 14963 29408
rect 14899 29348 14903 29404
rect 14903 29348 14959 29404
rect 14959 29348 14963 29404
rect 14899 29344 14963 29348
rect 13492 29140 13556 29204
rect 11652 29064 11716 29068
rect 11652 29008 11666 29064
rect 11666 29008 11716 29064
rect 11652 29004 11716 29008
rect 2665 28860 2729 28864
rect 2665 28804 2669 28860
rect 2669 28804 2725 28860
rect 2725 28804 2729 28860
rect 2665 28800 2729 28804
rect 2745 28860 2809 28864
rect 2745 28804 2749 28860
rect 2749 28804 2805 28860
rect 2805 28804 2809 28860
rect 2745 28800 2809 28804
rect 2825 28860 2889 28864
rect 2825 28804 2829 28860
rect 2829 28804 2885 28860
rect 2885 28804 2889 28860
rect 2825 28800 2889 28804
rect 2905 28860 2969 28864
rect 2905 28804 2909 28860
rect 2909 28804 2965 28860
rect 2965 28804 2969 28860
rect 2905 28800 2969 28804
rect 6092 28860 6156 28864
rect 6092 28804 6096 28860
rect 6096 28804 6152 28860
rect 6152 28804 6156 28860
rect 6092 28800 6156 28804
rect 6172 28860 6236 28864
rect 6172 28804 6176 28860
rect 6176 28804 6232 28860
rect 6232 28804 6236 28860
rect 6172 28800 6236 28804
rect 6252 28860 6316 28864
rect 6252 28804 6256 28860
rect 6256 28804 6312 28860
rect 6312 28804 6316 28860
rect 6252 28800 6316 28804
rect 6332 28860 6396 28864
rect 6332 28804 6336 28860
rect 6336 28804 6392 28860
rect 6392 28804 6396 28860
rect 6332 28800 6396 28804
rect 9519 28860 9583 28864
rect 9519 28804 9523 28860
rect 9523 28804 9579 28860
rect 9579 28804 9583 28860
rect 9519 28800 9583 28804
rect 9599 28860 9663 28864
rect 9599 28804 9603 28860
rect 9603 28804 9659 28860
rect 9659 28804 9663 28860
rect 9599 28800 9663 28804
rect 9679 28860 9743 28864
rect 9679 28804 9683 28860
rect 9683 28804 9739 28860
rect 9739 28804 9743 28860
rect 9679 28800 9743 28804
rect 9759 28860 9823 28864
rect 9759 28804 9763 28860
rect 9763 28804 9819 28860
rect 9819 28804 9823 28860
rect 9759 28800 9823 28804
rect 12946 28860 13010 28864
rect 12946 28804 12950 28860
rect 12950 28804 13006 28860
rect 13006 28804 13010 28860
rect 12946 28800 13010 28804
rect 13026 28860 13090 28864
rect 13026 28804 13030 28860
rect 13030 28804 13086 28860
rect 13086 28804 13090 28860
rect 13026 28800 13090 28804
rect 13106 28860 13170 28864
rect 13106 28804 13110 28860
rect 13110 28804 13166 28860
rect 13166 28804 13170 28860
rect 13106 28800 13170 28804
rect 13186 28860 13250 28864
rect 13186 28804 13190 28860
rect 13190 28804 13246 28860
rect 13246 28804 13250 28860
rect 13186 28800 13250 28804
rect 12756 28732 12820 28796
rect 1716 28460 1780 28524
rect 12756 28460 12820 28524
rect 4378 28316 4442 28320
rect 4378 28260 4382 28316
rect 4382 28260 4438 28316
rect 4438 28260 4442 28316
rect 4378 28256 4442 28260
rect 4458 28316 4522 28320
rect 4458 28260 4462 28316
rect 4462 28260 4518 28316
rect 4518 28260 4522 28316
rect 4458 28256 4522 28260
rect 4538 28316 4602 28320
rect 4538 28260 4542 28316
rect 4542 28260 4598 28316
rect 4598 28260 4602 28316
rect 4538 28256 4602 28260
rect 4618 28316 4682 28320
rect 4618 28260 4622 28316
rect 4622 28260 4678 28316
rect 4678 28260 4682 28316
rect 4618 28256 4682 28260
rect 7805 28316 7869 28320
rect 7805 28260 7809 28316
rect 7809 28260 7865 28316
rect 7865 28260 7869 28316
rect 7805 28256 7869 28260
rect 7885 28316 7949 28320
rect 7885 28260 7889 28316
rect 7889 28260 7945 28316
rect 7945 28260 7949 28316
rect 7885 28256 7949 28260
rect 7965 28316 8029 28320
rect 7965 28260 7969 28316
rect 7969 28260 8025 28316
rect 8025 28260 8029 28316
rect 7965 28256 8029 28260
rect 8045 28316 8109 28320
rect 8045 28260 8049 28316
rect 8049 28260 8105 28316
rect 8105 28260 8109 28316
rect 8045 28256 8109 28260
rect 11232 28316 11296 28320
rect 11232 28260 11236 28316
rect 11236 28260 11292 28316
rect 11292 28260 11296 28316
rect 11232 28256 11296 28260
rect 11312 28316 11376 28320
rect 11312 28260 11316 28316
rect 11316 28260 11372 28316
rect 11372 28260 11376 28316
rect 11312 28256 11376 28260
rect 11392 28316 11456 28320
rect 11392 28260 11396 28316
rect 11396 28260 11452 28316
rect 11452 28260 11456 28316
rect 11392 28256 11456 28260
rect 11472 28316 11536 28320
rect 11472 28260 11476 28316
rect 11476 28260 11532 28316
rect 11532 28260 11536 28316
rect 11472 28256 11536 28260
rect 14659 28316 14723 28320
rect 14659 28260 14663 28316
rect 14663 28260 14719 28316
rect 14719 28260 14723 28316
rect 14659 28256 14723 28260
rect 14739 28316 14803 28320
rect 14739 28260 14743 28316
rect 14743 28260 14799 28316
rect 14799 28260 14803 28316
rect 14739 28256 14803 28260
rect 14819 28316 14883 28320
rect 14819 28260 14823 28316
rect 14823 28260 14879 28316
rect 14879 28260 14883 28316
rect 14819 28256 14883 28260
rect 14899 28316 14963 28320
rect 14899 28260 14903 28316
rect 14903 28260 14959 28316
rect 14959 28260 14963 28316
rect 14899 28256 14963 28260
rect 13860 28188 13924 28252
rect 2665 27772 2729 27776
rect 2665 27716 2669 27772
rect 2669 27716 2725 27772
rect 2725 27716 2729 27772
rect 2665 27712 2729 27716
rect 2745 27772 2809 27776
rect 2745 27716 2749 27772
rect 2749 27716 2805 27772
rect 2805 27716 2809 27772
rect 2745 27712 2809 27716
rect 2825 27772 2889 27776
rect 2825 27716 2829 27772
rect 2829 27716 2885 27772
rect 2885 27716 2889 27772
rect 2825 27712 2889 27716
rect 2905 27772 2969 27776
rect 2905 27716 2909 27772
rect 2909 27716 2965 27772
rect 2965 27716 2969 27772
rect 2905 27712 2969 27716
rect 6092 27772 6156 27776
rect 6092 27716 6096 27772
rect 6096 27716 6152 27772
rect 6152 27716 6156 27772
rect 6092 27712 6156 27716
rect 6172 27772 6236 27776
rect 6172 27716 6176 27772
rect 6176 27716 6232 27772
rect 6232 27716 6236 27772
rect 6172 27712 6236 27716
rect 6252 27772 6316 27776
rect 6252 27716 6256 27772
rect 6256 27716 6312 27772
rect 6312 27716 6316 27772
rect 6252 27712 6316 27716
rect 6332 27772 6396 27776
rect 6332 27716 6336 27772
rect 6336 27716 6392 27772
rect 6392 27716 6396 27772
rect 6332 27712 6396 27716
rect 9519 27772 9583 27776
rect 9519 27716 9523 27772
rect 9523 27716 9579 27772
rect 9579 27716 9583 27772
rect 9519 27712 9583 27716
rect 9599 27772 9663 27776
rect 9599 27716 9603 27772
rect 9603 27716 9659 27772
rect 9659 27716 9663 27772
rect 9599 27712 9663 27716
rect 9679 27772 9743 27776
rect 9679 27716 9683 27772
rect 9683 27716 9739 27772
rect 9739 27716 9743 27772
rect 9679 27712 9743 27716
rect 9759 27772 9823 27776
rect 9759 27716 9763 27772
rect 9763 27716 9819 27772
rect 9819 27716 9823 27772
rect 9759 27712 9823 27716
rect 12946 27772 13010 27776
rect 12946 27716 12950 27772
rect 12950 27716 13006 27772
rect 13006 27716 13010 27772
rect 12946 27712 13010 27716
rect 13026 27772 13090 27776
rect 13026 27716 13030 27772
rect 13030 27716 13086 27772
rect 13086 27716 13090 27772
rect 13026 27712 13090 27716
rect 13106 27772 13170 27776
rect 13106 27716 13110 27772
rect 13110 27716 13166 27772
rect 13166 27716 13170 27772
rect 13106 27712 13170 27716
rect 13186 27772 13250 27776
rect 13186 27716 13190 27772
rect 13190 27716 13246 27772
rect 13246 27716 13250 27772
rect 13186 27712 13250 27716
rect 13676 27372 13740 27436
rect 4378 27228 4442 27232
rect 4378 27172 4382 27228
rect 4382 27172 4438 27228
rect 4438 27172 4442 27228
rect 4378 27168 4442 27172
rect 4458 27228 4522 27232
rect 4458 27172 4462 27228
rect 4462 27172 4518 27228
rect 4518 27172 4522 27228
rect 4458 27168 4522 27172
rect 4538 27228 4602 27232
rect 4538 27172 4542 27228
rect 4542 27172 4598 27228
rect 4598 27172 4602 27228
rect 4538 27168 4602 27172
rect 4618 27228 4682 27232
rect 4618 27172 4622 27228
rect 4622 27172 4678 27228
rect 4678 27172 4682 27228
rect 4618 27168 4682 27172
rect 7805 27228 7869 27232
rect 7805 27172 7809 27228
rect 7809 27172 7865 27228
rect 7865 27172 7869 27228
rect 7805 27168 7869 27172
rect 7885 27228 7949 27232
rect 7885 27172 7889 27228
rect 7889 27172 7945 27228
rect 7945 27172 7949 27228
rect 7885 27168 7949 27172
rect 7965 27228 8029 27232
rect 7965 27172 7969 27228
rect 7969 27172 8025 27228
rect 8025 27172 8029 27228
rect 7965 27168 8029 27172
rect 8045 27228 8109 27232
rect 8045 27172 8049 27228
rect 8049 27172 8105 27228
rect 8105 27172 8109 27228
rect 8045 27168 8109 27172
rect 11232 27228 11296 27232
rect 11232 27172 11236 27228
rect 11236 27172 11292 27228
rect 11292 27172 11296 27228
rect 11232 27168 11296 27172
rect 11312 27228 11376 27232
rect 11312 27172 11316 27228
rect 11316 27172 11372 27228
rect 11372 27172 11376 27228
rect 11312 27168 11376 27172
rect 11392 27228 11456 27232
rect 11392 27172 11396 27228
rect 11396 27172 11452 27228
rect 11452 27172 11456 27228
rect 11392 27168 11456 27172
rect 11472 27228 11536 27232
rect 11472 27172 11476 27228
rect 11476 27172 11532 27228
rect 11532 27172 11536 27228
rect 11472 27168 11536 27172
rect 14659 27228 14723 27232
rect 14659 27172 14663 27228
rect 14663 27172 14719 27228
rect 14719 27172 14723 27228
rect 14659 27168 14723 27172
rect 14739 27228 14803 27232
rect 14739 27172 14743 27228
rect 14743 27172 14799 27228
rect 14799 27172 14803 27228
rect 14739 27168 14803 27172
rect 14819 27228 14883 27232
rect 14819 27172 14823 27228
rect 14823 27172 14879 27228
rect 14879 27172 14883 27228
rect 14819 27168 14883 27172
rect 14899 27228 14963 27232
rect 14899 27172 14903 27228
rect 14903 27172 14959 27228
rect 14959 27172 14963 27228
rect 14899 27168 14963 27172
rect 2665 26684 2729 26688
rect 2665 26628 2669 26684
rect 2669 26628 2725 26684
rect 2725 26628 2729 26684
rect 2665 26624 2729 26628
rect 2745 26684 2809 26688
rect 2745 26628 2749 26684
rect 2749 26628 2805 26684
rect 2805 26628 2809 26684
rect 2745 26624 2809 26628
rect 2825 26684 2889 26688
rect 2825 26628 2829 26684
rect 2829 26628 2885 26684
rect 2885 26628 2889 26684
rect 2825 26624 2889 26628
rect 2905 26684 2969 26688
rect 2905 26628 2909 26684
rect 2909 26628 2965 26684
rect 2965 26628 2969 26684
rect 2905 26624 2969 26628
rect 6092 26684 6156 26688
rect 6092 26628 6096 26684
rect 6096 26628 6152 26684
rect 6152 26628 6156 26684
rect 6092 26624 6156 26628
rect 6172 26684 6236 26688
rect 6172 26628 6176 26684
rect 6176 26628 6232 26684
rect 6232 26628 6236 26684
rect 6172 26624 6236 26628
rect 6252 26684 6316 26688
rect 6252 26628 6256 26684
rect 6256 26628 6312 26684
rect 6312 26628 6316 26684
rect 6252 26624 6316 26628
rect 6332 26684 6396 26688
rect 6332 26628 6336 26684
rect 6336 26628 6392 26684
rect 6392 26628 6396 26684
rect 6332 26624 6396 26628
rect 9519 26684 9583 26688
rect 9519 26628 9523 26684
rect 9523 26628 9579 26684
rect 9579 26628 9583 26684
rect 9519 26624 9583 26628
rect 9599 26684 9663 26688
rect 9599 26628 9603 26684
rect 9603 26628 9659 26684
rect 9659 26628 9663 26684
rect 9599 26624 9663 26628
rect 9679 26684 9743 26688
rect 9679 26628 9683 26684
rect 9683 26628 9739 26684
rect 9739 26628 9743 26684
rect 9679 26624 9743 26628
rect 9759 26684 9823 26688
rect 9759 26628 9763 26684
rect 9763 26628 9819 26684
rect 9819 26628 9823 26684
rect 9759 26624 9823 26628
rect 12946 26684 13010 26688
rect 12946 26628 12950 26684
rect 12950 26628 13006 26684
rect 13006 26628 13010 26684
rect 12946 26624 13010 26628
rect 13026 26684 13090 26688
rect 13026 26628 13030 26684
rect 13030 26628 13086 26684
rect 13086 26628 13090 26684
rect 13026 26624 13090 26628
rect 13106 26684 13170 26688
rect 13106 26628 13110 26684
rect 13110 26628 13166 26684
rect 13166 26628 13170 26684
rect 13106 26624 13170 26628
rect 13186 26684 13250 26688
rect 13186 26628 13190 26684
rect 13190 26628 13246 26684
rect 13246 26628 13250 26684
rect 13186 26624 13250 26628
rect 3924 26284 3988 26348
rect 4378 26140 4442 26144
rect 4378 26084 4382 26140
rect 4382 26084 4438 26140
rect 4438 26084 4442 26140
rect 4378 26080 4442 26084
rect 4458 26140 4522 26144
rect 4458 26084 4462 26140
rect 4462 26084 4518 26140
rect 4518 26084 4522 26140
rect 4458 26080 4522 26084
rect 4538 26140 4602 26144
rect 4538 26084 4542 26140
rect 4542 26084 4598 26140
rect 4598 26084 4602 26140
rect 4538 26080 4602 26084
rect 4618 26140 4682 26144
rect 4618 26084 4622 26140
rect 4622 26084 4678 26140
rect 4678 26084 4682 26140
rect 4618 26080 4682 26084
rect 7805 26140 7869 26144
rect 7805 26084 7809 26140
rect 7809 26084 7865 26140
rect 7865 26084 7869 26140
rect 7805 26080 7869 26084
rect 7885 26140 7949 26144
rect 7885 26084 7889 26140
rect 7889 26084 7945 26140
rect 7945 26084 7949 26140
rect 7885 26080 7949 26084
rect 7965 26140 8029 26144
rect 7965 26084 7969 26140
rect 7969 26084 8025 26140
rect 8025 26084 8029 26140
rect 7965 26080 8029 26084
rect 8045 26140 8109 26144
rect 8045 26084 8049 26140
rect 8049 26084 8105 26140
rect 8105 26084 8109 26140
rect 8045 26080 8109 26084
rect 11232 26140 11296 26144
rect 11232 26084 11236 26140
rect 11236 26084 11292 26140
rect 11292 26084 11296 26140
rect 11232 26080 11296 26084
rect 11312 26140 11376 26144
rect 11312 26084 11316 26140
rect 11316 26084 11372 26140
rect 11372 26084 11376 26140
rect 11312 26080 11376 26084
rect 11392 26140 11456 26144
rect 11392 26084 11396 26140
rect 11396 26084 11452 26140
rect 11452 26084 11456 26140
rect 11392 26080 11456 26084
rect 11472 26140 11536 26144
rect 11472 26084 11476 26140
rect 11476 26084 11532 26140
rect 11532 26084 11536 26140
rect 11472 26080 11536 26084
rect 14659 26140 14723 26144
rect 14659 26084 14663 26140
rect 14663 26084 14719 26140
rect 14719 26084 14723 26140
rect 14659 26080 14723 26084
rect 14739 26140 14803 26144
rect 14739 26084 14743 26140
rect 14743 26084 14799 26140
rect 14799 26084 14803 26140
rect 14739 26080 14803 26084
rect 14819 26140 14883 26144
rect 14819 26084 14823 26140
rect 14823 26084 14879 26140
rect 14879 26084 14883 26140
rect 14819 26080 14883 26084
rect 14899 26140 14963 26144
rect 14899 26084 14903 26140
rect 14903 26084 14959 26140
rect 14959 26084 14963 26140
rect 14899 26080 14963 26084
rect 2665 25596 2729 25600
rect 2665 25540 2669 25596
rect 2669 25540 2725 25596
rect 2725 25540 2729 25596
rect 2665 25536 2729 25540
rect 2745 25596 2809 25600
rect 2745 25540 2749 25596
rect 2749 25540 2805 25596
rect 2805 25540 2809 25596
rect 2745 25536 2809 25540
rect 2825 25596 2889 25600
rect 2825 25540 2829 25596
rect 2829 25540 2885 25596
rect 2885 25540 2889 25596
rect 2825 25536 2889 25540
rect 2905 25596 2969 25600
rect 2905 25540 2909 25596
rect 2909 25540 2965 25596
rect 2965 25540 2969 25596
rect 2905 25536 2969 25540
rect 6092 25596 6156 25600
rect 6092 25540 6096 25596
rect 6096 25540 6152 25596
rect 6152 25540 6156 25596
rect 6092 25536 6156 25540
rect 6172 25596 6236 25600
rect 6172 25540 6176 25596
rect 6176 25540 6232 25596
rect 6232 25540 6236 25596
rect 6172 25536 6236 25540
rect 6252 25596 6316 25600
rect 6252 25540 6256 25596
rect 6256 25540 6312 25596
rect 6312 25540 6316 25596
rect 6252 25536 6316 25540
rect 6332 25596 6396 25600
rect 6332 25540 6336 25596
rect 6336 25540 6392 25596
rect 6392 25540 6396 25596
rect 6332 25536 6396 25540
rect 9519 25596 9583 25600
rect 9519 25540 9523 25596
rect 9523 25540 9579 25596
rect 9579 25540 9583 25596
rect 9519 25536 9583 25540
rect 9599 25596 9663 25600
rect 9599 25540 9603 25596
rect 9603 25540 9659 25596
rect 9659 25540 9663 25596
rect 9599 25536 9663 25540
rect 9679 25596 9743 25600
rect 9679 25540 9683 25596
rect 9683 25540 9739 25596
rect 9739 25540 9743 25596
rect 9679 25536 9743 25540
rect 9759 25596 9823 25600
rect 9759 25540 9763 25596
rect 9763 25540 9819 25596
rect 9819 25540 9823 25596
rect 9759 25536 9823 25540
rect 12946 25596 13010 25600
rect 12946 25540 12950 25596
rect 12950 25540 13006 25596
rect 13006 25540 13010 25596
rect 12946 25536 13010 25540
rect 13026 25596 13090 25600
rect 13026 25540 13030 25596
rect 13030 25540 13086 25596
rect 13086 25540 13090 25596
rect 13026 25536 13090 25540
rect 13106 25596 13170 25600
rect 13106 25540 13110 25596
rect 13110 25540 13166 25596
rect 13166 25540 13170 25596
rect 13106 25536 13170 25540
rect 13186 25596 13250 25600
rect 13186 25540 13190 25596
rect 13190 25540 13246 25596
rect 13246 25540 13250 25596
rect 13186 25536 13250 25540
rect 6500 25196 6564 25260
rect 10548 25060 10612 25124
rect 4378 25052 4442 25056
rect 4378 24996 4382 25052
rect 4382 24996 4438 25052
rect 4438 24996 4442 25052
rect 4378 24992 4442 24996
rect 4458 25052 4522 25056
rect 4458 24996 4462 25052
rect 4462 24996 4518 25052
rect 4518 24996 4522 25052
rect 4458 24992 4522 24996
rect 4538 25052 4602 25056
rect 4538 24996 4542 25052
rect 4542 24996 4598 25052
rect 4598 24996 4602 25052
rect 4538 24992 4602 24996
rect 4618 25052 4682 25056
rect 4618 24996 4622 25052
rect 4622 24996 4678 25052
rect 4678 24996 4682 25052
rect 4618 24992 4682 24996
rect 7805 25052 7869 25056
rect 7805 24996 7809 25052
rect 7809 24996 7865 25052
rect 7865 24996 7869 25052
rect 7805 24992 7869 24996
rect 7885 25052 7949 25056
rect 7885 24996 7889 25052
rect 7889 24996 7945 25052
rect 7945 24996 7949 25052
rect 7885 24992 7949 24996
rect 7965 25052 8029 25056
rect 7965 24996 7969 25052
rect 7969 24996 8025 25052
rect 8025 24996 8029 25052
rect 7965 24992 8029 24996
rect 8045 25052 8109 25056
rect 8045 24996 8049 25052
rect 8049 24996 8105 25052
rect 8105 24996 8109 25052
rect 8045 24992 8109 24996
rect 11232 25052 11296 25056
rect 11232 24996 11236 25052
rect 11236 24996 11292 25052
rect 11292 24996 11296 25052
rect 11232 24992 11296 24996
rect 11312 25052 11376 25056
rect 11312 24996 11316 25052
rect 11316 24996 11372 25052
rect 11372 24996 11376 25052
rect 11312 24992 11376 24996
rect 11392 25052 11456 25056
rect 11392 24996 11396 25052
rect 11396 24996 11452 25052
rect 11452 24996 11456 25052
rect 11392 24992 11456 24996
rect 11472 25052 11536 25056
rect 11472 24996 11476 25052
rect 11476 24996 11532 25052
rect 11532 24996 11536 25052
rect 11472 24992 11536 24996
rect 14659 25052 14723 25056
rect 14659 24996 14663 25052
rect 14663 24996 14719 25052
rect 14719 24996 14723 25052
rect 14659 24992 14723 24996
rect 14739 25052 14803 25056
rect 14739 24996 14743 25052
rect 14743 24996 14799 25052
rect 14799 24996 14803 25052
rect 14739 24992 14803 24996
rect 14819 25052 14883 25056
rect 14819 24996 14823 25052
rect 14823 24996 14879 25052
rect 14879 24996 14883 25052
rect 14819 24992 14883 24996
rect 14899 25052 14963 25056
rect 14899 24996 14903 25052
rect 14903 24996 14959 25052
rect 14959 24996 14963 25052
rect 14899 24992 14963 24996
rect 10548 24652 10612 24716
rect 13492 24652 13556 24716
rect 2665 24508 2729 24512
rect 2665 24452 2669 24508
rect 2669 24452 2725 24508
rect 2725 24452 2729 24508
rect 2665 24448 2729 24452
rect 2745 24508 2809 24512
rect 2745 24452 2749 24508
rect 2749 24452 2805 24508
rect 2805 24452 2809 24508
rect 2745 24448 2809 24452
rect 2825 24508 2889 24512
rect 2825 24452 2829 24508
rect 2829 24452 2885 24508
rect 2885 24452 2889 24508
rect 2825 24448 2889 24452
rect 2905 24508 2969 24512
rect 2905 24452 2909 24508
rect 2909 24452 2965 24508
rect 2965 24452 2969 24508
rect 2905 24448 2969 24452
rect 6092 24508 6156 24512
rect 6092 24452 6096 24508
rect 6096 24452 6152 24508
rect 6152 24452 6156 24508
rect 6092 24448 6156 24452
rect 6172 24508 6236 24512
rect 6172 24452 6176 24508
rect 6176 24452 6232 24508
rect 6232 24452 6236 24508
rect 6172 24448 6236 24452
rect 6252 24508 6316 24512
rect 6252 24452 6256 24508
rect 6256 24452 6312 24508
rect 6312 24452 6316 24508
rect 6252 24448 6316 24452
rect 6332 24508 6396 24512
rect 6332 24452 6336 24508
rect 6336 24452 6392 24508
rect 6392 24452 6396 24508
rect 6332 24448 6396 24452
rect 9519 24508 9583 24512
rect 9519 24452 9523 24508
rect 9523 24452 9579 24508
rect 9579 24452 9583 24508
rect 9519 24448 9583 24452
rect 9599 24508 9663 24512
rect 9599 24452 9603 24508
rect 9603 24452 9659 24508
rect 9659 24452 9663 24508
rect 9599 24448 9663 24452
rect 9679 24508 9743 24512
rect 9679 24452 9683 24508
rect 9683 24452 9739 24508
rect 9739 24452 9743 24508
rect 9679 24448 9743 24452
rect 9759 24508 9823 24512
rect 9759 24452 9763 24508
rect 9763 24452 9819 24508
rect 9819 24452 9823 24508
rect 9759 24448 9823 24452
rect 12946 24508 13010 24512
rect 12946 24452 12950 24508
rect 12950 24452 13006 24508
rect 13006 24452 13010 24508
rect 12946 24448 13010 24452
rect 13026 24508 13090 24512
rect 13026 24452 13030 24508
rect 13030 24452 13086 24508
rect 13086 24452 13090 24508
rect 13026 24448 13090 24452
rect 13106 24508 13170 24512
rect 13106 24452 13110 24508
rect 13110 24452 13166 24508
rect 13166 24452 13170 24508
rect 13106 24448 13170 24452
rect 13186 24508 13250 24512
rect 13186 24452 13190 24508
rect 13190 24452 13246 24508
rect 13246 24452 13250 24508
rect 13186 24448 13250 24452
rect 7420 23972 7484 24036
rect 4378 23964 4442 23968
rect 4378 23908 4382 23964
rect 4382 23908 4438 23964
rect 4438 23908 4442 23964
rect 4378 23904 4442 23908
rect 4458 23964 4522 23968
rect 4458 23908 4462 23964
rect 4462 23908 4518 23964
rect 4518 23908 4522 23964
rect 4458 23904 4522 23908
rect 4538 23964 4602 23968
rect 4538 23908 4542 23964
rect 4542 23908 4598 23964
rect 4598 23908 4602 23964
rect 4538 23904 4602 23908
rect 4618 23964 4682 23968
rect 4618 23908 4622 23964
rect 4622 23908 4678 23964
rect 4678 23908 4682 23964
rect 4618 23904 4682 23908
rect 7805 23964 7869 23968
rect 7805 23908 7809 23964
rect 7809 23908 7865 23964
rect 7865 23908 7869 23964
rect 7805 23904 7869 23908
rect 7885 23964 7949 23968
rect 7885 23908 7889 23964
rect 7889 23908 7945 23964
rect 7945 23908 7949 23964
rect 7885 23904 7949 23908
rect 7965 23964 8029 23968
rect 7965 23908 7969 23964
rect 7969 23908 8025 23964
rect 8025 23908 8029 23964
rect 7965 23904 8029 23908
rect 8045 23964 8109 23968
rect 8045 23908 8049 23964
rect 8049 23908 8105 23964
rect 8105 23908 8109 23964
rect 8045 23904 8109 23908
rect 11232 23964 11296 23968
rect 11232 23908 11236 23964
rect 11236 23908 11292 23964
rect 11292 23908 11296 23964
rect 11232 23904 11296 23908
rect 11312 23964 11376 23968
rect 11312 23908 11316 23964
rect 11316 23908 11372 23964
rect 11372 23908 11376 23964
rect 11312 23904 11376 23908
rect 11392 23964 11456 23968
rect 11392 23908 11396 23964
rect 11396 23908 11452 23964
rect 11452 23908 11456 23964
rect 11392 23904 11456 23908
rect 11472 23964 11536 23968
rect 11472 23908 11476 23964
rect 11476 23908 11532 23964
rect 11532 23908 11536 23964
rect 11472 23904 11536 23908
rect 7420 23836 7484 23900
rect 14659 23964 14723 23968
rect 14659 23908 14663 23964
rect 14663 23908 14719 23964
rect 14719 23908 14723 23964
rect 14659 23904 14723 23908
rect 14739 23964 14803 23968
rect 14739 23908 14743 23964
rect 14743 23908 14799 23964
rect 14799 23908 14803 23964
rect 14739 23904 14803 23908
rect 14819 23964 14883 23968
rect 14819 23908 14823 23964
rect 14823 23908 14879 23964
rect 14879 23908 14883 23964
rect 14819 23904 14883 23908
rect 14899 23964 14963 23968
rect 14899 23908 14903 23964
rect 14903 23908 14959 23964
rect 14959 23908 14963 23964
rect 14899 23904 14963 23908
rect 2665 23420 2729 23424
rect 2665 23364 2669 23420
rect 2669 23364 2725 23420
rect 2725 23364 2729 23420
rect 2665 23360 2729 23364
rect 2745 23420 2809 23424
rect 2745 23364 2749 23420
rect 2749 23364 2805 23420
rect 2805 23364 2809 23420
rect 2745 23360 2809 23364
rect 2825 23420 2889 23424
rect 2825 23364 2829 23420
rect 2829 23364 2885 23420
rect 2885 23364 2889 23420
rect 2825 23360 2889 23364
rect 2905 23420 2969 23424
rect 2905 23364 2909 23420
rect 2909 23364 2965 23420
rect 2965 23364 2969 23420
rect 2905 23360 2969 23364
rect 6092 23420 6156 23424
rect 6092 23364 6096 23420
rect 6096 23364 6152 23420
rect 6152 23364 6156 23420
rect 6092 23360 6156 23364
rect 6172 23420 6236 23424
rect 6172 23364 6176 23420
rect 6176 23364 6232 23420
rect 6232 23364 6236 23420
rect 6172 23360 6236 23364
rect 6252 23420 6316 23424
rect 6252 23364 6256 23420
rect 6256 23364 6312 23420
rect 6312 23364 6316 23420
rect 6252 23360 6316 23364
rect 6332 23420 6396 23424
rect 6332 23364 6336 23420
rect 6336 23364 6392 23420
rect 6392 23364 6396 23420
rect 6332 23360 6396 23364
rect 9519 23420 9583 23424
rect 9519 23364 9523 23420
rect 9523 23364 9579 23420
rect 9579 23364 9583 23420
rect 9519 23360 9583 23364
rect 9599 23420 9663 23424
rect 9599 23364 9603 23420
rect 9603 23364 9659 23420
rect 9659 23364 9663 23420
rect 9599 23360 9663 23364
rect 9679 23420 9743 23424
rect 9679 23364 9683 23420
rect 9683 23364 9739 23420
rect 9739 23364 9743 23420
rect 9679 23360 9743 23364
rect 9759 23420 9823 23424
rect 9759 23364 9763 23420
rect 9763 23364 9819 23420
rect 9819 23364 9823 23420
rect 9759 23360 9823 23364
rect 12946 23420 13010 23424
rect 12946 23364 12950 23420
rect 12950 23364 13006 23420
rect 13006 23364 13010 23420
rect 12946 23360 13010 23364
rect 13026 23420 13090 23424
rect 13026 23364 13030 23420
rect 13030 23364 13086 23420
rect 13086 23364 13090 23420
rect 13026 23360 13090 23364
rect 13106 23420 13170 23424
rect 13106 23364 13110 23420
rect 13110 23364 13166 23420
rect 13166 23364 13170 23420
rect 13106 23360 13170 23364
rect 13186 23420 13250 23424
rect 13186 23364 13190 23420
rect 13190 23364 13246 23420
rect 13246 23364 13250 23420
rect 13186 23360 13250 23364
rect 7236 23156 7300 23220
rect 8892 23080 8956 23084
rect 8892 23024 8906 23080
rect 8906 23024 8956 23080
rect 8892 23020 8956 23024
rect 11652 23020 11716 23084
rect 12572 23080 12636 23084
rect 12572 23024 12622 23080
rect 12622 23024 12636 23080
rect 12572 23020 12636 23024
rect 4378 22876 4442 22880
rect 4378 22820 4382 22876
rect 4382 22820 4438 22876
rect 4438 22820 4442 22876
rect 4378 22816 4442 22820
rect 4458 22876 4522 22880
rect 4458 22820 4462 22876
rect 4462 22820 4518 22876
rect 4518 22820 4522 22876
rect 4458 22816 4522 22820
rect 4538 22876 4602 22880
rect 4538 22820 4542 22876
rect 4542 22820 4598 22876
rect 4598 22820 4602 22876
rect 4538 22816 4602 22820
rect 4618 22876 4682 22880
rect 4618 22820 4622 22876
rect 4622 22820 4678 22876
rect 4678 22820 4682 22876
rect 4618 22816 4682 22820
rect 7805 22876 7869 22880
rect 7805 22820 7809 22876
rect 7809 22820 7865 22876
rect 7865 22820 7869 22876
rect 7805 22816 7869 22820
rect 7885 22876 7949 22880
rect 7885 22820 7889 22876
rect 7889 22820 7945 22876
rect 7945 22820 7949 22876
rect 7885 22816 7949 22820
rect 7965 22876 8029 22880
rect 7965 22820 7969 22876
rect 7969 22820 8025 22876
rect 8025 22820 8029 22876
rect 7965 22816 8029 22820
rect 8045 22876 8109 22880
rect 8045 22820 8049 22876
rect 8049 22820 8105 22876
rect 8105 22820 8109 22876
rect 8045 22816 8109 22820
rect 11232 22876 11296 22880
rect 11232 22820 11236 22876
rect 11236 22820 11292 22876
rect 11292 22820 11296 22876
rect 11232 22816 11296 22820
rect 11312 22876 11376 22880
rect 11312 22820 11316 22876
rect 11316 22820 11372 22876
rect 11372 22820 11376 22876
rect 11312 22816 11376 22820
rect 11392 22876 11456 22880
rect 11392 22820 11396 22876
rect 11396 22820 11452 22876
rect 11452 22820 11456 22876
rect 11392 22816 11456 22820
rect 11472 22876 11536 22880
rect 11472 22820 11476 22876
rect 11476 22820 11532 22876
rect 11532 22820 11536 22876
rect 11472 22816 11536 22820
rect 14659 22876 14723 22880
rect 14659 22820 14663 22876
rect 14663 22820 14719 22876
rect 14719 22820 14723 22876
rect 14659 22816 14723 22820
rect 14739 22876 14803 22880
rect 14739 22820 14743 22876
rect 14743 22820 14799 22876
rect 14799 22820 14803 22876
rect 14739 22816 14803 22820
rect 14819 22876 14883 22880
rect 14819 22820 14823 22876
rect 14823 22820 14879 22876
rect 14879 22820 14883 22876
rect 14819 22816 14883 22820
rect 14899 22876 14963 22880
rect 14899 22820 14903 22876
rect 14903 22820 14959 22876
rect 14959 22820 14963 22876
rect 14899 22816 14963 22820
rect 9260 22612 9324 22676
rect 11836 22612 11900 22676
rect 8892 22476 8956 22540
rect 2665 22332 2729 22336
rect 2665 22276 2669 22332
rect 2669 22276 2725 22332
rect 2725 22276 2729 22332
rect 2665 22272 2729 22276
rect 2745 22332 2809 22336
rect 2745 22276 2749 22332
rect 2749 22276 2805 22332
rect 2805 22276 2809 22332
rect 2745 22272 2809 22276
rect 2825 22332 2889 22336
rect 2825 22276 2829 22332
rect 2829 22276 2885 22332
rect 2885 22276 2889 22332
rect 2825 22272 2889 22276
rect 2905 22332 2969 22336
rect 2905 22276 2909 22332
rect 2909 22276 2965 22332
rect 2965 22276 2969 22332
rect 2905 22272 2969 22276
rect 6092 22332 6156 22336
rect 6092 22276 6096 22332
rect 6096 22276 6152 22332
rect 6152 22276 6156 22332
rect 6092 22272 6156 22276
rect 6172 22332 6236 22336
rect 6172 22276 6176 22332
rect 6176 22276 6232 22332
rect 6232 22276 6236 22332
rect 6172 22272 6236 22276
rect 6252 22332 6316 22336
rect 6252 22276 6256 22332
rect 6256 22276 6312 22332
rect 6312 22276 6316 22332
rect 6252 22272 6316 22276
rect 6332 22332 6396 22336
rect 6332 22276 6336 22332
rect 6336 22276 6392 22332
rect 6392 22276 6396 22332
rect 6332 22272 6396 22276
rect 9519 22332 9583 22336
rect 9519 22276 9523 22332
rect 9523 22276 9579 22332
rect 9579 22276 9583 22332
rect 9519 22272 9583 22276
rect 9599 22332 9663 22336
rect 9599 22276 9603 22332
rect 9603 22276 9659 22332
rect 9659 22276 9663 22332
rect 9599 22272 9663 22276
rect 9679 22332 9743 22336
rect 9679 22276 9683 22332
rect 9683 22276 9739 22332
rect 9739 22276 9743 22332
rect 9679 22272 9743 22276
rect 9759 22332 9823 22336
rect 9759 22276 9763 22332
rect 9763 22276 9819 22332
rect 9819 22276 9823 22332
rect 9759 22272 9823 22276
rect 12946 22332 13010 22336
rect 12946 22276 12950 22332
rect 12950 22276 13006 22332
rect 13006 22276 13010 22332
rect 12946 22272 13010 22276
rect 13026 22332 13090 22336
rect 13026 22276 13030 22332
rect 13030 22276 13086 22332
rect 13086 22276 13090 22332
rect 13026 22272 13090 22276
rect 13106 22332 13170 22336
rect 13106 22276 13110 22332
rect 13110 22276 13166 22332
rect 13166 22276 13170 22332
rect 13106 22272 13170 22276
rect 13186 22332 13250 22336
rect 13186 22276 13190 22332
rect 13190 22276 13246 22332
rect 13246 22276 13250 22332
rect 13186 22272 13250 22276
rect 12756 22068 12820 22132
rect 7604 21992 7668 21996
rect 7604 21936 7618 21992
rect 7618 21936 7668 21992
rect 7604 21932 7668 21936
rect 4378 21788 4442 21792
rect 4378 21732 4382 21788
rect 4382 21732 4438 21788
rect 4438 21732 4442 21788
rect 4378 21728 4442 21732
rect 4458 21788 4522 21792
rect 4458 21732 4462 21788
rect 4462 21732 4518 21788
rect 4518 21732 4522 21788
rect 4458 21728 4522 21732
rect 4538 21788 4602 21792
rect 4538 21732 4542 21788
rect 4542 21732 4598 21788
rect 4598 21732 4602 21788
rect 4538 21728 4602 21732
rect 4618 21788 4682 21792
rect 4618 21732 4622 21788
rect 4622 21732 4678 21788
rect 4678 21732 4682 21788
rect 4618 21728 4682 21732
rect 7805 21788 7869 21792
rect 7805 21732 7809 21788
rect 7809 21732 7865 21788
rect 7865 21732 7869 21788
rect 7805 21728 7869 21732
rect 7885 21788 7949 21792
rect 7885 21732 7889 21788
rect 7889 21732 7945 21788
rect 7945 21732 7949 21788
rect 7885 21728 7949 21732
rect 7965 21788 8029 21792
rect 7965 21732 7969 21788
rect 7969 21732 8025 21788
rect 8025 21732 8029 21788
rect 7965 21728 8029 21732
rect 8045 21788 8109 21792
rect 8045 21732 8049 21788
rect 8049 21732 8105 21788
rect 8105 21732 8109 21788
rect 8045 21728 8109 21732
rect 11232 21788 11296 21792
rect 11232 21732 11236 21788
rect 11236 21732 11292 21788
rect 11292 21732 11296 21788
rect 11232 21728 11296 21732
rect 11312 21788 11376 21792
rect 11312 21732 11316 21788
rect 11316 21732 11372 21788
rect 11372 21732 11376 21788
rect 11312 21728 11376 21732
rect 11392 21788 11456 21792
rect 11392 21732 11396 21788
rect 11396 21732 11452 21788
rect 11452 21732 11456 21788
rect 11392 21728 11456 21732
rect 11472 21788 11536 21792
rect 11472 21732 11476 21788
rect 11476 21732 11532 21788
rect 11532 21732 11536 21788
rect 11472 21728 11536 21732
rect 14659 21788 14723 21792
rect 14659 21732 14663 21788
rect 14663 21732 14719 21788
rect 14719 21732 14723 21788
rect 14659 21728 14723 21732
rect 14739 21788 14803 21792
rect 14739 21732 14743 21788
rect 14743 21732 14799 21788
rect 14799 21732 14803 21788
rect 14739 21728 14803 21732
rect 14819 21788 14883 21792
rect 14819 21732 14823 21788
rect 14823 21732 14879 21788
rect 14879 21732 14883 21788
rect 14819 21728 14883 21732
rect 14899 21788 14963 21792
rect 14899 21732 14903 21788
rect 14903 21732 14959 21788
rect 14959 21732 14963 21788
rect 14899 21728 14963 21732
rect 9996 21660 10060 21724
rect 2665 21244 2729 21248
rect 2665 21188 2669 21244
rect 2669 21188 2725 21244
rect 2725 21188 2729 21244
rect 2665 21184 2729 21188
rect 2745 21244 2809 21248
rect 2745 21188 2749 21244
rect 2749 21188 2805 21244
rect 2805 21188 2809 21244
rect 2745 21184 2809 21188
rect 2825 21244 2889 21248
rect 2825 21188 2829 21244
rect 2829 21188 2885 21244
rect 2885 21188 2889 21244
rect 2825 21184 2889 21188
rect 2905 21244 2969 21248
rect 2905 21188 2909 21244
rect 2909 21188 2965 21244
rect 2965 21188 2969 21244
rect 2905 21184 2969 21188
rect 6092 21244 6156 21248
rect 6092 21188 6096 21244
rect 6096 21188 6152 21244
rect 6152 21188 6156 21244
rect 6092 21184 6156 21188
rect 6172 21244 6236 21248
rect 6172 21188 6176 21244
rect 6176 21188 6232 21244
rect 6232 21188 6236 21244
rect 6172 21184 6236 21188
rect 6252 21244 6316 21248
rect 6252 21188 6256 21244
rect 6256 21188 6312 21244
rect 6312 21188 6316 21244
rect 6252 21184 6316 21188
rect 6332 21244 6396 21248
rect 6332 21188 6336 21244
rect 6336 21188 6392 21244
rect 6392 21188 6396 21244
rect 6332 21184 6396 21188
rect 9519 21244 9583 21248
rect 9519 21188 9523 21244
rect 9523 21188 9579 21244
rect 9579 21188 9583 21244
rect 9519 21184 9583 21188
rect 9599 21244 9663 21248
rect 9599 21188 9603 21244
rect 9603 21188 9659 21244
rect 9659 21188 9663 21244
rect 9599 21184 9663 21188
rect 9679 21244 9743 21248
rect 9679 21188 9683 21244
rect 9683 21188 9739 21244
rect 9739 21188 9743 21244
rect 9679 21184 9743 21188
rect 9759 21244 9823 21248
rect 9759 21188 9763 21244
rect 9763 21188 9819 21244
rect 9819 21188 9823 21244
rect 9759 21184 9823 21188
rect 12946 21244 13010 21248
rect 12946 21188 12950 21244
rect 12950 21188 13006 21244
rect 13006 21188 13010 21244
rect 12946 21184 13010 21188
rect 13026 21244 13090 21248
rect 13026 21188 13030 21244
rect 13030 21188 13086 21244
rect 13086 21188 13090 21244
rect 13026 21184 13090 21188
rect 13106 21244 13170 21248
rect 13106 21188 13110 21244
rect 13110 21188 13166 21244
rect 13166 21188 13170 21244
rect 13106 21184 13170 21188
rect 13186 21244 13250 21248
rect 13186 21188 13190 21244
rect 13190 21188 13246 21244
rect 13246 21188 13250 21244
rect 13186 21184 13250 21188
rect 12204 21176 12268 21180
rect 12204 21120 12254 21176
rect 12254 21120 12268 21176
rect 12204 21116 12268 21120
rect 4378 20700 4442 20704
rect 4378 20644 4382 20700
rect 4382 20644 4438 20700
rect 4438 20644 4442 20700
rect 4378 20640 4442 20644
rect 4458 20700 4522 20704
rect 4458 20644 4462 20700
rect 4462 20644 4518 20700
rect 4518 20644 4522 20700
rect 4458 20640 4522 20644
rect 4538 20700 4602 20704
rect 4538 20644 4542 20700
rect 4542 20644 4598 20700
rect 4598 20644 4602 20700
rect 4538 20640 4602 20644
rect 4618 20700 4682 20704
rect 4618 20644 4622 20700
rect 4622 20644 4678 20700
rect 4678 20644 4682 20700
rect 4618 20640 4682 20644
rect 7805 20700 7869 20704
rect 7805 20644 7809 20700
rect 7809 20644 7865 20700
rect 7865 20644 7869 20700
rect 7805 20640 7869 20644
rect 7885 20700 7949 20704
rect 7885 20644 7889 20700
rect 7889 20644 7945 20700
rect 7945 20644 7949 20700
rect 7885 20640 7949 20644
rect 7965 20700 8029 20704
rect 7965 20644 7969 20700
rect 7969 20644 8025 20700
rect 8025 20644 8029 20700
rect 7965 20640 8029 20644
rect 8045 20700 8109 20704
rect 8045 20644 8049 20700
rect 8049 20644 8105 20700
rect 8105 20644 8109 20700
rect 8045 20640 8109 20644
rect 11232 20700 11296 20704
rect 11232 20644 11236 20700
rect 11236 20644 11292 20700
rect 11292 20644 11296 20700
rect 11232 20640 11296 20644
rect 11312 20700 11376 20704
rect 11312 20644 11316 20700
rect 11316 20644 11372 20700
rect 11372 20644 11376 20700
rect 11312 20640 11376 20644
rect 11392 20700 11456 20704
rect 11392 20644 11396 20700
rect 11396 20644 11452 20700
rect 11452 20644 11456 20700
rect 11392 20640 11456 20644
rect 11472 20700 11536 20704
rect 11472 20644 11476 20700
rect 11476 20644 11532 20700
rect 11532 20644 11536 20700
rect 11472 20640 11536 20644
rect 14659 20700 14723 20704
rect 14659 20644 14663 20700
rect 14663 20644 14719 20700
rect 14719 20644 14723 20700
rect 14659 20640 14723 20644
rect 14739 20700 14803 20704
rect 14739 20644 14743 20700
rect 14743 20644 14799 20700
rect 14799 20644 14803 20700
rect 14739 20640 14803 20644
rect 14819 20700 14883 20704
rect 14819 20644 14823 20700
rect 14823 20644 14879 20700
rect 14879 20644 14883 20700
rect 14819 20640 14883 20644
rect 14899 20700 14963 20704
rect 14899 20644 14903 20700
rect 14903 20644 14959 20700
rect 14959 20644 14963 20700
rect 14899 20640 14963 20644
rect 2665 20156 2729 20160
rect 2665 20100 2669 20156
rect 2669 20100 2725 20156
rect 2725 20100 2729 20156
rect 2665 20096 2729 20100
rect 2745 20156 2809 20160
rect 2745 20100 2749 20156
rect 2749 20100 2805 20156
rect 2805 20100 2809 20156
rect 2745 20096 2809 20100
rect 2825 20156 2889 20160
rect 2825 20100 2829 20156
rect 2829 20100 2885 20156
rect 2885 20100 2889 20156
rect 2825 20096 2889 20100
rect 2905 20156 2969 20160
rect 2905 20100 2909 20156
rect 2909 20100 2965 20156
rect 2965 20100 2969 20156
rect 2905 20096 2969 20100
rect 6092 20156 6156 20160
rect 6092 20100 6096 20156
rect 6096 20100 6152 20156
rect 6152 20100 6156 20156
rect 6092 20096 6156 20100
rect 6172 20156 6236 20160
rect 6172 20100 6176 20156
rect 6176 20100 6232 20156
rect 6232 20100 6236 20156
rect 6172 20096 6236 20100
rect 6252 20156 6316 20160
rect 6252 20100 6256 20156
rect 6256 20100 6312 20156
rect 6312 20100 6316 20156
rect 6252 20096 6316 20100
rect 6332 20156 6396 20160
rect 6332 20100 6336 20156
rect 6336 20100 6392 20156
rect 6392 20100 6396 20156
rect 6332 20096 6396 20100
rect 9519 20156 9583 20160
rect 9519 20100 9523 20156
rect 9523 20100 9579 20156
rect 9579 20100 9583 20156
rect 9519 20096 9583 20100
rect 9599 20156 9663 20160
rect 9599 20100 9603 20156
rect 9603 20100 9659 20156
rect 9659 20100 9663 20156
rect 9599 20096 9663 20100
rect 9679 20156 9743 20160
rect 9679 20100 9683 20156
rect 9683 20100 9739 20156
rect 9739 20100 9743 20156
rect 9679 20096 9743 20100
rect 9759 20156 9823 20160
rect 9759 20100 9763 20156
rect 9763 20100 9819 20156
rect 9819 20100 9823 20156
rect 9759 20096 9823 20100
rect 12946 20156 13010 20160
rect 12946 20100 12950 20156
rect 12950 20100 13006 20156
rect 13006 20100 13010 20156
rect 12946 20096 13010 20100
rect 13026 20156 13090 20160
rect 13026 20100 13030 20156
rect 13030 20100 13086 20156
rect 13086 20100 13090 20156
rect 13026 20096 13090 20100
rect 13106 20156 13170 20160
rect 13106 20100 13110 20156
rect 13110 20100 13166 20156
rect 13166 20100 13170 20156
rect 13106 20096 13170 20100
rect 13186 20156 13250 20160
rect 13186 20100 13190 20156
rect 13190 20100 13246 20156
rect 13246 20100 13250 20156
rect 13186 20096 13250 20100
rect 13676 19892 13740 19956
rect 4378 19612 4442 19616
rect 4378 19556 4382 19612
rect 4382 19556 4438 19612
rect 4438 19556 4442 19612
rect 4378 19552 4442 19556
rect 4458 19612 4522 19616
rect 4458 19556 4462 19612
rect 4462 19556 4518 19612
rect 4518 19556 4522 19612
rect 4458 19552 4522 19556
rect 4538 19612 4602 19616
rect 4538 19556 4542 19612
rect 4542 19556 4598 19612
rect 4598 19556 4602 19612
rect 4538 19552 4602 19556
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 7805 19612 7869 19616
rect 7805 19556 7809 19612
rect 7809 19556 7865 19612
rect 7865 19556 7869 19612
rect 7805 19552 7869 19556
rect 7885 19612 7949 19616
rect 7885 19556 7889 19612
rect 7889 19556 7945 19612
rect 7945 19556 7949 19612
rect 7885 19552 7949 19556
rect 7965 19612 8029 19616
rect 7965 19556 7969 19612
rect 7969 19556 8025 19612
rect 8025 19556 8029 19612
rect 7965 19552 8029 19556
rect 8045 19612 8109 19616
rect 8045 19556 8049 19612
rect 8049 19556 8105 19612
rect 8105 19556 8109 19612
rect 8045 19552 8109 19556
rect 11232 19612 11296 19616
rect 11232 19556 11236 19612
rect 11236 19556 11292 19612
rect 11292 19556 11296 19612
rect 11232 19552 11296 19556
rect 11312 19612 11376 19616
rect 11312 19556 11316 19612
rect 11316 19556 11372 19612
rect 11372 19556 11376 19612
rect 11312 19552 11376 19556
rect 11392 19612 11456 19616
rect 11392 19556 11396 19612
rect 11396 19556 11452 19612
rect 11452 19556 11456 19612
rect 11392 19552 11456 19556
rect 11472 19612 11536 19616
rect 11472 19556 11476 19612
rect 11476 19556 11532 19612
rect 11532 19556 11536 19612
rect 11472 19552 11536 19556
rect 14659 19612 14723 19616
rect 14659 19556 14663 19612
rect 14663 19556 14719 19612
rect 14719 19556 14723 19612
rect 14659 19552 14723 19556
rect 14739 19612 14803 19616
rect 14739 19556 14743 19612
rect 14743 19556 14799 19612
rect 14799 19556 14803 19612
rect 14739 19552 14803 19556
rect 14819 19612 14883 19616
rect 14819 19556 14823 19612
rect 14823 19556 14879 19612
rect 14879 19556 14883 19612
rect 14819 19552 14883 19556
rect 14899 19612 14963 19616
rect 14899 19556 14903 19612
rect 14903 19556 14959 19612
rect 14959 19556 14963 19612
rect 14899 19552 14963 19556
rect 9076 19544 9140 19548
rect 9076 19488 9090 19544
rect 9090 19488 9140 19544
rect 9076 19484 9140 19488
rect 9996 19544 10060 19548
rect 9996 19488 10046 19544
rect 10046 19488 10060 19544
rect 9996 19484 10060 19488
rect 2665 19068 2729 19072
rect 2665 19012 2669 19068
rect 2669 19012 2725 19068
rect 2725 19012 2729 19068
rect 2665 19008 2729 19012
rect 2745 19068 2809 19072
rect 2745 19012 2749 19068
rect 2749 19012 2805 19068
rect 2805 19012 2809 19068
rect 2745 19008 2809 19012
rect 2825 19068 2889 19072
rect 2825 19012 2829 19068
rect 2829 19012 2885 19068
rect 2885 19012 2889 19068
rect 2825 19008 2889 19012
rect 2905 19068 2969 19072
rect 2905 19012 2909 19068
rect 2909 19012 2965 19068
rect 2965 19012 2969 19068
rect 2905 19008 2969 19012
rect 6092 19068 6156 19072
rect 6092 19012 6096 19068
rect 6096 19012 6152 19068
rect 6152 19012 6156 19068
rect 6092 19008 6156 19012
rect 6172 19068 6236 19072
rect 6172 19012 6176 19068
rect 6176 19012 6232 19068
rect 6232 19012 6236 19068
rect 6172 19008 6236 19012
rect 6252 19068 6316 19072
rect 6252 19012 6256 19068
rect 6256 19012 6312 19068
rect 6312 19012 6316 19068
rect 6252 19008 6316 19012
rect 6332 19068 6396 19072
rect 6332 19012 6336 19068
rect 6336 19012 6392 19068
rect 6392 19012 6396 19068
rect 6332 19008 6396 19012
rect 9519 19068 9583 19072
rect 9519 19012 9523 19068
rect 9523 19012 9579 19068
rect 9579 19012 9583 19068
rect 9519 19008 9583 19012
rect 9599 19068 9663 19072
rect 9599 19012 9603 19068
rect 9603 19012 9659 19068
rect 9659 19012 9663 19068
rect 9599 19008 9663 19012
rect 9679 19068 9743 19072
rect 9679 19012 9683 19068
rect 9683 19012 9739 19068
rect 9739 19012 9743 19068
rect 9679 19008 9743 19012
rect 9759 19068 9823 19072
rect 9759 19012 9763 19068
rect 9763 19012 9819 19068
rect 9819 19012 9823 19068
rect 9759 19008 9823 19012
rect 12946 19068 13010 19072
rect 12946 19012 12950 19068
rect 12950 19012 13006 19068
rect 13006 19012 13010 19068
rect 12946 19008 13010 19012
rect 13026 19068 13090 19072
rect 13026 19012 13030 19068
rect 13030 19012 13086 19068
rect 13086 19012 13090 19068
rect 13026 19008 13090 19012
rect 13106 19068 13170 19072
rect 13106 19012 13110 19068
rect 13110 19012 13166 19068
rect 13166 19012 13170 19068
rect 13106 19008 13170 19012
rect 13186 19068 13250 19072
rect 13186 19012 13190 19068
rect 13190 19012 13246 19068
rect 13246 19012 13250 19068
rect 13186 19008 13250 19012
rect 11836 18940 11900 19004
rect 7420 18864 7484 18868
rect 7420 18808 7434 18864
rect 7434 18808 7484 18864
rect 7420 18804 7484 18808
rect 12572 18804 12636 18868
rect 7420 18668 7484 18732
rect 10732 18668 10796 18732
rect 4378 18524 4442 18528
rect 4378 18468 4382 18524
rect 4382 18468 4438 18524
rect 4438 18468 4442 18524
rect 4378 18464 4442 18468
rect 4458 18524 4522 18528
rect 4458 18468 4462 18524
rect 4462 18468 4518 18524
rect 4518 18468 4522 18524
rect 4458 18464 4522 18468
rect 4538 18524 4602 18528
rect 4538 18468 4542 18524
rect 4542 18468 4598 18524
rect 4598 18468 4602 18524
rect 4538 18464 4602 18468
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 7805 18524 7869 18528
rect 7805 18468 7809 18524
rect 7809 18468 7865 18524
rect 7865 18468 7869 18524
rect 7805 18464 7869 18468
rect 7885 18524 7949 18528
rect 7885 18468 7889 18524
rect 7889 18468 7945 18524
rect 7945 18468 7949 18524
rect 7885 18464 7949 18468
rect 7965 18524 8029 18528
rect 7965 18468 7969 18524
rect 7969 18468 8025 18524
rect 8025 18468 8029 18524
rect 7965 18464 8029 18468
rect 8045 18524 8109 18528
rect 8045 18468 8049 18524
rect 8049 18468 8105 18524
rect 8105 18468 8109 18524
rect 8045 18464 8109 18468
rect 11232 18524 11296 18528
rect 11232 18468 11236 18524
rect 11236 18468 11292 18524
rect 11292 18468 11296 18524
rect 11232 18464 11296 18468
rect 11312 18524 11376 18528
rect 11312 18468 11316 18524
rect 11316 18468 11372 18524
rect 11372 18468 11376 18524
rect 11312 18464 11376 18468
rect 11392 18524 11456 18528
rect 11392 18468 11396 18524
rect 11396 18468 11452 18524
rect 11452 18468 11456 18524
rect 11392 18464 11456 18468
rect 11472 18524 11536 18528
rect 11472 18468 11476 18524
rect 11476 18468 11532 18524
rect 11532 18468 11536 18524
rect 11472 18464 11536 18468
rect 14659 18524 14723 18528
rect 14659 18468 14663 18524
rect 14663 18468 14719 18524
rect 14719 18468 14723 18524
rect 14659 18464 14723 18468
rect 14739 18524 14803 18528
rect 14739 18468 14743 18524
rect 14743 18468 14799 18524
rect 14799 18468 14803 18524
rect 14739 18464 14803 18468
rect 14819 18524 14883 18528
rect 14819 18468 14823 18524
rect 14823 18468 14879 18524
rect 14879 18468 14883 18524
rect 14819 18464 14883 18468
rect 14899 18524 14963 18528
rect 14899 18468 14903 18524
rect 14903 18468 14959 18524
rect 14959 18468 14963 18524
rect 14899 18464 14963 18468
rect 2665 17980 2729 17984
rect 2665 17924 2669 17980
rect 2669 17924 2725 17980
rect 2725 17924 2729 17980
rect 2665 17920 2729 17924
rect 2745 17980 2809 17984
rect 2745 17924 2749 17980
rect 2749 17924 2805 17980
rect 2805 17924 2809 17980
rect 2745 17920 2809 17924
rect 2825 17980 2889 17984
rect 2825 17924 2829 17980
rect 2829 17924 2885 17980
rect 2885 17924 2889 17980
rect 2825 17920 2889 17924
rect 2905 17980 2969 17984
rect 2905 17924 2909 17980
rect 2909 17924 2965 17980
rect 2965 17924 2969 17980
rect 2905 17920 2969 17924
rect 6092 17980 6156 17984
rect 6092 17924 6096 17980
rect 6096 17924 6152 17980
rect 6152 17924 6156 17980
rect 6092 17920 6156 17924
rect 6172 17980 6236 17984
rect 6172 17924 6176 17980
rect 6176 17924 6232 17980
rect 6232 17924 6236 17980
rect 6172 17920 6236 17924
rect 6252 17980 6316 17984
rect 6252 17924 6256 17980
rect 6256 17924 6312 17980
rect 6312 17924 6316 17980
rect 6252 17920 6316 17924
rect 6332 17980 6396 17984
rect 6332 17924 6336 17980
rect 6336 17924 6392 17980
rect 6392 17924 6396 17980
rect 6332 17920 6396 17924
rect 9519 17980 9583 17984
rect 9519 17924 9523 17980
rect 9523 17924 9579 17980
rect 9579 17924 9583 17980
rect 9519 17920 9583 17924
rect 9599 17980 9663 17984
rect 9599 17924 9603 17980
rect 9603 17924 9659 17980
rect 9659 17924 9663 17980
rect 9599 17920 9663 17924
rect 9679 17980 9743 17984
rect 9679 17924 9683 17980
rect 9683 17924 9739 17980
rect 9739 17924 9743 17980
rect 9679 17920 9743 17924
rect 9759 17980 9823 17984
rect 9759 17924 9763 17980
rect 9763 17924 9819 17980
rect 9819 17924 9823 17980
rect 9759 17920 9823 17924
rect 12946 17980 13010 17984
rect 12946 17924 12950 17980
rect 12950 17924 13006 17980
rect 13006 17924 13010 17980
rect 12946 17920 13010 17924
rect 13026 17980 13090 17984
rect 13026 17924 13030 17980
rect 13030 17924 13086 17980
rect 13086 17924 13090 17980
rect 13026 17920 13090 17924
rect 13106 17980 13170 17984
rect 13106 17924 13110 17980
rect 13110 17924 13166 17980
rect 13166 17924 13170 17980
rect 13106 17920 13170 17924
rect 13186 17980 13250 17984
rect 13186 17924 13190 17980
rect 13190 17924 13246 17980
rect 13246 17924 13250 17980
rect 13186 17920 13250 17924
rect 13860 17912 13924 17916
rect 13860 17856 13874 17912
rect 13874 17856 13924 17912
rect 13860 17852 13924 17856
rect 6500 17640 6564 17644
rect 10548 17716 10612 17780
rect 6500 17584 6514 17640
rect 6514 17584 6564 17640
rect 6500 17580 6564 17584
rect 11836 17580 11900 17644
rect 14228 17504 14292 17508
rect 14228 17448 14242 17504
rect 14242 17448 14292 17504
rect 14228 17444 14292 17448
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 13492 17308 13556 17372
rect 11652 17036 11716 17100
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 12204 16764 12268 16828
rect 14044 16628 14108 16692
rect 7604 16552 7668 16556
rect 7604 16496 7618 16552
rect 7618 16496 7668 16552
rect 7604 16492 7668 16496
rect 9260 16552 9324 16556
rect 9260 16496 9274 16552
rect 9274 16496 9324 16552
rect 9260 16492 9324 16496
rect 10548 16356 10612 16420
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 12756 15268 12820 15332
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 8892 15132 8956 15196
rect 12756 15132 12820 15196
rect 13676 14860 13740 14924
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 10732 14316 10796 14380
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 10548 13772 10612 13836
rect 14228 13832 14292 13836
rect 14228 13776 14242 13832
rect 14242 13776 14292 13832
rect 14228 13772 14292 13776
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 7420 12820 7484 12884
rect 3924 12684 3988 12748
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 14044 12140 14108 12204
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 13676 11928 13740 11932
rect 13676 11872 13726 11928
rect 13726 11872 13740 11928
rect 13676 11868 13740 11872
rect 13492 11732 13556 11796
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 2268 10644 2332 10708
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 12756 10024 12820 10028
rect 12756 9968 12806 10024
rect 12806 9968 12820 10024
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 11652 9692 11716 9756
rect 1716 9616 1780 9620
rect 1716 9560 1766 9616
rect 1766 9560 1780 9616
rect 1716 9556 1780 9560
rect 12756 9964 12820 9968
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 11652 9284 11716 9348
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12204 9012 12268 9076
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 12204 8604 12268 8668
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 6684 3436 6748 3500
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 10916 2620 10980 2684
rect 11836 2680 11900 2684
rect 11836 2624 11850 2680
rect 11850 2624 11900 2680
rect 11836 2620 11900 2624
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
rect 2665 1660 2729 1664
rect 2665 1604 2669 1660
rect 2669 1604 2725 1660
rect 2725 1604 2729 1660
rect 2665 1600 2729 1604
rect 2745 1660 2809 1664
rect 2745 1604 2749 1660
rect 2749 1604 2805 1660
rect 2805 1604 2809 1660
rect 2745 1600 2809 1604
rect 2825 1660 2889 1664
rect 2825 1604 2829 1660
rect 2829 1604 2885 1660
rect 2885 1604 2889 1660
rect 2825 1600 2889 1604
rect 2905 1660 2969 1664
rect 2905 1604 2909 1660
rect 2909 1604 2965 1660
rect 2965 1604 2969 1660
rect 2905 1600 2969 1604
rect 6092 1660 6156 1664
rect 6092 1604 6096 1660
rect 6096 1604 6152 1660
rect 6152 1604 6156 1660
rect 6092 1600 6156 1604
rect 6172 1660 6236 1664
rect 6172 1604 6176 1660
rect 6176 1604 6232 1660
rect 6232 1604 6236 1660
rect 6172 1600 6236 1604
rect 6252 1660 6316 1664
rect 6252 1604 6256 1660
rect 6256 1604 6312 1660
rect 6312 1604 6316 1660
rect 6252 1600 6316 1604
rect 6332 1660 6396 1664
rect 6332 1604 6336 1660
rect 6336 1604 6392 1660
rect 6392 1604 6396 1660
rect 6332 1600 6396 1604
rect 9519 1660 9583 1664
rect 9519 1604 9523 1660
rect 9523 1604 9579 1660
rect 9579 1604 9583 1660
rect 9519 1600 9583 1604
rect 9599 1660 9663 1664
rect 9599 1604 9603 1660
rect 9603 1604 9659 1660
rect 9659 1604 9663 1660
rect 9599 1600 9663 1604
rect 9679 1660 9743 1664
rect 9679 1604 9683 1660
rect 9683 1604 9739 1660
rect 9739 1604 9743 1660
rect 9679 1600 9743 1604
rect 9759 1660 9823 1664
rect 9759 1604 9763 1660
rect 9763 1604 9819 1660
rect 9819 1604 9823 1660
rect 9759 1600 9823 1604
rect 12946 1660 13010 1664
rect 12946 1604 12950 1660
rect 12950 1604 13006 1660
rect 13006 1604 13010 1660
rect 12946 1600 13010 1604
rect 13026 1660 13090 1664
rect 13026 1604 13030 1660
rect 13030 1604 13086 1660
rect 13086 1604 13090 1660
rect 13026 1600 13090 1604
rect 13106 1660 13170 1664
rect 13106 1604 13110 1660
rect 13110 1604 13166 1660
rect 13166 1604 13170 1660
rect 13106 1600 13170 1604
rect 13186 1660 13250 1664
rect 13186 1604 13190 1660
rect 13190 1604 13246 1660
rect 13246 1604 13250 1660
rect 13186 1600 13250 1604
rect 4844 1260 4908 1324
rect 5396 1320 5460 1324
rect 5396 1264 5410 1320
rect 5410 1264 5460 1320
rect 5396 1260 5460 1264
rect 4378 1116 4442 1120
rect 4378 1060 4382 1116
rect 4382 1060 4438 1116
rect 4438 1060 4442 1116
rect 4378 1056 4442 1060
rect 4458 1116 4522 1120
rect 4458 1060 4462 1116
rect 4462 1060 4518 1116
rect 4518 1060 4522 1116
rect 4458 1056 4522 1060
rect 4538 1116 4602 1120
rect 4538 1060 4542 1116
rect 4542 1060 4598 1116
rect 4598 1060 4602 1116
rect 4538 1056 4602 1060
rect 4618 1116 4682 1120
rect 4618 1060 4622 1116
rect 4622 1060 4678 1116
rect 4678 1060 4682 1116
rect 4618 1056 4682 1060
rect 7805 1116 7869 1120
rect 7805 1060 7809 1116
rect 7809 1060 7865 1116
rect 7865 1060 7869 1116
rect 7805 1056 7869 1060
rect 7885 1116 7949 1120
rect 7885 1060 7889 1116
rect 7889 1060 7945 1116
rect 7945 1060 7949 1116
rect 7885 1056 7949 1060
rect 7965 1116 8029 1120
rect 7965 1060 7969 1116
rect 7969 1060 8025 1116
rect 8025 1060 8029 1116
rect 7965 1056 8029 1060
rect 8045 1116 8109 1120
rect 8045 1060 8049 1116
rect 8049 1060 8105 1116
rect 8105 1060 8109 1116
rect 8045 1056 8109 1060
rect 11232 1116 11296 1120
rect 11232 1060 11236 1116
rect 11236 1060 11292 1116
rect 11292 1060 11296 1116
rect 11232 1056 11296 1060
rect 11312 1116 11376 1120
rect 11312 1060 11316 1116
rect 11316 1060 11372 1116
rect 11372 1060 11376 1116
rect 11312 1056 11376 1060
rect 11392 1116 11456 1120
rect 11392 1060 11396 1116
rect 11396 1060 11452 1116
rect 11452 1060 11456 1116
rect 11392 1056 11456 1060
rect 11472 1116 11536 1120
rect 11472 1060 11476 1116
rect 11476 1060 11532 1116
rect 11532 1060 11536 1116
rect 11472 1056 11536 1060
rect 14659 1116 14723 1120
rect 14659 1060 14663 1116
rect 14663 1060 14719 1116
rect 14719 1060 14723 1116
rect 14659 1056 14723 1060
rect 14739 1116 14803 1120
rect 14739 1060 14743 1116
rect 14743 1060 14799 1116
rect 14799 1060 14803 1116
rect 14739 1056 14803 1060
rect 14819 1116 14883 1120
rect 14819 1060 14823 1116
rect 14823 1060 14879 1116
rect 14879 1060 14883 1116
rect 14819 1056 14883 1060
rect 14899 1116 14963 1120
rect 14899 1060 14903 1116
rect 14903 1060 14959 1116
rect 14959 1060 14963 1116
rect 14899 1056 14963 1060
<< metal4 >>
rect 2657 43008 2977 43568
rect 2657 42944 2665 43008
rect 2729 42944 2745 43008
rect 2809 42944 2825 43008
rect 2889 42944 2905 43008
rect 2969 42944 2977 43008
rect 2657 41920 2977 42944
rect 2657 41856 2665 41920
rect 2729 41856 2745 41920
rect 2809 41856 2825 41920
rect 2889 41856 2905 41920
rect 2969 41856 2977 41920
rect 2267 41716 2333 41717
rect 2267 41652 2268 41716
rect 2332 41652 2333 41716
rect 2267 41651 2333 41652
rect 1715 28524 1781 28525
rect 1715 28460 1716 28524
rect 1780 28460 1781 28524
rect 1715 28459 1781 28460
rect 1718 9621 1778 28459
rect 2270 10709 2330 41651
rect 2657 40832 2977 41856
rect 2657 40768 2665 40832
rect 2729 40768 2745 40832
rect 2809 40768 2825 40832
rect 2889 40768 2905 40832
rect 2969 40768 2977 40832
rect 2657 39744 2977 40768
rect 2657 39680 2665 39744
rect 2729 39680 2745 39744
rect 2809 39680 2825 39744
rect 2889 39680 2905 39744
rect 2969 39680 2977 39744
rect 2657 38656 2977 39680
rect 2657 38592 2665 38656
rect 2729 38592 2745 38656
rect 2809 38592 2825 38656
rect 2889 38592 2905 38656
rect 2969 38592 2977 38656
rect 2657 37568 2977 38592
rect 2657 37504 2665 37568
rect 2729 37504 2745 37568
rect 2809 37504 2825 37568
rect 2889 37504 2905 37568
rect 2969 37504 2977 37568
rect 2657 36480 2977 37504
rect 2657 36416 2665 36480
rect 2729 36416 2745 36480
rect 2809 36416 2825 36480
rect 2889 36416 2905 36480
rect 2969 36416 2977 36480
rect 2657 35392 2977 36416
rect 2657 35328 2665 35392
rect 2729 35328 2745 35392
rect 2809 35328 2825 35392
rect 2889 35328 2905 35392
rect 2969 35328 2977 35392
rect 2657 34304 2977 35328
rect 2657 34240 2665 34304
rect 2729 34240 2745 34304
rect 2809 34240 2825 34304
rect 2889 34240 2905 34304
rect 2969 34240 2977 34304
rect 2657 33216 2977 34240
rect 2657 33152 2665 33216
rect 2729 33152 2745 33216
rect 2809 33152 2825 33216
rect 2889 33152 2905 33216
rect 2969 33152 2977 33216
rect 2657 32128 2977 33152
rect 2657 32064 2665 32128
rect 2729 32064 2745 32128
rect 2809 32064 2825 32128
rect 2889 32064 2905 32128
rect 2969 32064 2977 32128
rect 2657 31040 2977 32064
rect 2657 30976 2665 31040
rect 2729 30976 2745 31040
rect 2809 30976 2825 31040
rect 2889 30976 2905 31040
rect 2969 30976 2977 31040
rect 2657 29952 2977 30976
rect 2657 29888 2665 29952
rect 2729 29888 2745 29952
rect 2809 29888 2825 29952
rect 2889 29888 2905 29952
rect 2969 29888 2977 29952
rect 2657 28864 2977 29888
rect 2657 28800 2665 28864
rect 2729 28800 2745 28864
rect 2809 28800 2825 28864
rect 2889 28800 2905 28864
rect 2969 28800 2977 28864
rect 2657 27776 2977 28800
rect 2657 27712 2665 27776
rect 2729 27712 2745 27776
rect 2809 27712 2825 27776
rect 2889 27712 2905 27776
rect 2969 27712 2977 27776
rect 2657 26688 2977 27712
rect 2657 26624 2665 26688
rect 2729 26624 2745 26688
rect 2809 26624 2825 26688
rect 2889 26624 2905 26688
rect 2969 26624 2977 26688
rect 2657 25600 2977 26624
rect 4370 43552 4690 43568
rect 4370 43488 4378 43552
rect 4442 43488 4458 43552
rect 4522 43488 4538 43552
rect 4602 43488 4618 43552
rect 4682 43488 4690 43552
rect 4370 42464 4690 43488
rect 4370 42400 4378 42464
rect 4442 42400 4458 42464
rect 4522 42400 4538 42464
rect 4602 42400 4618 42464
rect 4682 42400 4690 42464
rect 4370 41376 4690 42400
rect 6084 43008 6404 43568
rect 6084 42944 6092 43008
rect 6156 42944 6172 43008
rect 6236 42944 6252 43008
rect 6316 42944 6332 43008
rect 6396 42944 6404 43008
rect 6084 41920 6404 42944
rect 7797 43552 8117 43568
rect 7797 43488 7805 43552
rect 7869 43488 7885 43552
rect 7949 43488 7965 43552
rect 8029 43488 8045 43552
rect 8109 43488 8117 43552
rect 6683 42668 6749 42669
rect 6683 42604 6684 42668
rect 6748 42604 6749 42668
rect 6683 42603 6749 42604
rect 6084 41856 6092 41920
rect 6156 41856 6172 41920
rect 6236 41856 6252 41920
rect 6316 41856 6332 41920
rect 6396 41856 6404 41920
rect 4843 41580 4909 41581
rect 4843 41516 4844 41580
rect 4908 41516 4909 41580
rect 4843 41515 4909 41516
rect 4370 41312 4378 41376
rect 4442 41312 4458 41376
rect 4522 41312 4538 41376
rect 4602 41312 4618 41376
rect 4682 41312 4690 41376
rect 4370 40288 4690 41312
rect 4370 40224 4378 40288
rect 4442 40224 4458 40288
rect 4522 40224 4538 40288
rect 4602 40224 4618 40288
rect 4682 40224 4690 40288
rect 4370 39200 4690 40224
rect 4370 39136 4378 39200
rect 4442 39136 4458 39200
rect 4522 39136 4538 39200
rect 4602 39136 4618 39200
rect 4682 39136 4690 39200
rect 4370 38112 4690 39136
rect 4370 38048 4378 38112
rect 4442 38048 4458 38112
rect 4522 38048 4538 38112
rect 4602 38048 4618 38112
rect 4682 38048 4690 38112
rect 4370 37024 4690 38048
rect 4370 36960 4378 37024
rect 4442 36960 4458 37024
rect 4522 36960 4538 37024
rect 4602 36960 4618 37024
rect 4682 36960 4690 37024
rect 4370 35936 4690 36960
rect 4370 35872 4378 35936
rect 4442 35872 4458 35936
rect 4522 35872 4538 35936
rect 4602 35872 4618 35936
rect 4682 35872 4690 35936
rect 4370 34848 4690 35872
rect 4370 34784 4378 34848
rect 4442 34784 4458 34848
rect 4522 34784 4538 34848
rect 4602 34784 4618 34848
rect 4682 34784 4690 34848
rect 4370 33760 4690 34784
rect 4370 33696 4378 33760
rect 4442 33696 4458 33760
rect 4522 33696 4538 33760
rect 4602 33696 4618 33760
rect 4682 33696 4690 33760
rect 4370 32672 4690 33696
rect 4370 32608 4378 32672
rect 4442 32608 4458 32672
rect 4522 32608 4538 32672
rect 4602 32608 4618 32672
rect 4682 32608 4690 32672
rect 4370 31584 4690 32608
rect 4370 31520 4378 31584
rect 4442 31520 4458 31584
rect 4522 31520 4538 31584
rect 4602 31520 4618 31584
rect 4682 31520 4690 31584
rect 4370 30496 4690 31520
rect 4370 30432 4378 30496
rect 4442 30432 4458 30496
rect 4522 30432 4538 30496
rect 4602 30432 4618 30496
rect 4682 30432 4690 30496
rect 4370 29408 4690 30432
rect 4370 29344 4378 29408
rect 4442 29344 4458 29408
rect 4522 29344 4538 29408
rect 4602 29344 4618 29408
rect 4682 29344 4690 29408
rect 4370 28320 4690 29344
rect 4370 28256 4378 28320
rect 4442 28256 4458 28320
rect 4522 28256 4538 28320
rect 4602 28256 4618 28320
rect 4682 28256 4690 28320
rect 4370 27232 4690 28256
rect 4370 27168 4378 27232
rect 4442 27168 4458 27232
rect 4522 27168 4538 27232
rect 4602 27168 4618 27232
rect 4682 27168 4690 27232
rect 3923 26348 3989 26349
rect 3923 26284 3924 26348
rect 3988 26284 3989 26348
rect 3923 26283 3989 26284
rect 2657 25536 2665 25600
rect 2729 25536 2745 25600
rect 2809 25536 2825 25600
rect 2889 25536 2905 25600
rect 2969 25536 2977 25600
rect 2657 24512 2977 25536
rect 2657 24448 2665 24512
rect 2729 24448 2745 24512
rect 2809 24448 2825 24512
rect 2889 24448 2905 24512
rect 2969 24448 2977 24512
rect 2657 23424 2977 24448
rect 2657 23360 2665 23424
rect 2729 23360 2745 23424
rect 2809 23360 2825 23424
rect 2889 23360 2905 23424
rect 2969 23360 2977 23424
rect 2657 22336 2977 23360
rect 2657 22272 2665 22336
rect 2729 22272 2745 22336
rect 2809 22272 2825 22336
rect 2889 22272 2905 22336
rect 2969 22272 2977 22336
rect 2657 21248 2977 22272
rect 2657 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2977 21248
rect 2657 20160 2977 21184
rect 2657 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2977 20160
rect 2657 19072 2977 20096
rect 2657 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2977 19072
rect 2657 17984 2977 19008
rect 2657 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2977 17984
rect 2657 16896 2977 17920
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 2657 13632 2977 14656
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 3926 12749 3986 26283
rect 4370 26144 4690 27168
rect 4370 26080 4378 26144
rect 4442 26080 4458 26144
rect 4522 26080 4538 26144
rect 4602 26080 4618 26144
rect 4682 26080 4690 26144
rect 4370 25056 4690 26080
rect 4370 24992 4378 25056
rect 4442 24992 4458 25056
rect 4522 24992 4538 25056
rect 4602 24992 4618 25056
rect 4682 24992 4690 25056
rect 4370 23968 4690 24992
rect 4370 23904 4378 23968
rect 4442 23904 4458 23968
rect 4522 23904 4538 23968
rect 4602 23904 4618 23968
rect 4682 23904 4690 23968
rect 4370 22880 4690 23904
rect 4370 22816 4378 22880
rect 4442 22816 4458 22880
rect 4522 22816 4538 22880
rect 4602 22816 4618 22880
rect 4682 22816 4690 22880
rect 4370 21792 4690 22816
rect 4370 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4690 21792
rect 4370 20704 4690 21728
rect 4370 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4690 20704
rect 4370 19616 4690 20640
rect 4370 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4690 19616
rect 4370 18528 4690 19552
rect 4370 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4690 18528
rect 4370 17440 4690 18464
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 3923 12748 3989 12749
rect 3923 12684 3924 12748
rect 3988 12684 3989 12748
rect 3923 12683 3989 12684
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2267 10708 2333 10709
rect 2267 10644 2268 10708
rect 2332 10644 2333 10708
rect 2267 10643 2333 10644
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 1715 9620 1781 9621
rect 1715 9556 1716 9620
rect 1780 9556 1781 9620
rect 1715 9555 1781 9556
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 1664 2977 2688
rect 2657 1600 2665 1664
rect 2729 1600 2745 1664
rect 2809 1600 2825 1664
rect 2889 1600 2905 1664
rect 2969 1600 2977 1664
rect 2657 1040 2977 1600
rect 4370 12000 4690 13024
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 1120 4690 2144
rect 4846 1325 4906 41515
rect 5395 41444 5461 41445
rect 5395 41380 5396 41444
rect 5460 41380 5461 41444
rect 5395 41379 5461 41380
rect 5398 1325 5458 41379
rect 6084 40832 6404 41856
rect 6084 40768 6092 40832
rect 6156 40768 6172 40832
rect 6236 40768 6252 40832
rect 6316 40768 6332 40832
rect 6396 40768 6404 40832
rect 6084 39744 6404 40768
rect 6084 39680 6092 39744
rect 6156 39680 6172 39744
rect 6236 39680 6252 39744
rect 6316 39680 6332 39744
rect 6396 39680 6404 39744
rect 6084 38656 6404 39680
rect 6084 38592 6092 38656
rect 6156 38592 6172 38656
rect 6236 38592 6252 38656
rect 6316 38592 6332 38656
rect 6396 38592 6404 38656
rect 6084 37568 6404 38592
rect 6084 37504 6092 37568
rect 6156 37504 6172 37568
rect 6236 37504 6252 37568
rect 6316 37504 6332 37568
rect 6396 37504 6404 37568
rect 6084 36480 6404 37504
rect 6084 36416 6092 36480
rect 6156 36416 6172 36480
rect 6236 36416 6252 36480
rect 6316 36416 6332 36480
rect 6396 36416 6404 36480
rect 6084 35392 6404 36416
rect 6084 35328 6092 35392
rect 6156 35328 6172 35392
rect 6236 35328 6252 35392
rect 6316 35328 6332 35392
rect 6396 35328 6404 35392
rect 6084 34304 6404 35328
rect 6084 34240 6092 34304
rect 6156 34240 6172 34304
rect 6236 34240 6252 34304
rect 6316 34240 6332 34304
rect 6396 34240 6404 34304
rect 6084 33216 6404 34240
rect 6084 33152 6092 33216
rect 6156 33152 6172 33216
rect 6236 33152 6252 33216
rect 6316 33152 6332 33216
rect 6396 33152 6404 33216
rect 6084 32128 6404 33152
rect 6084 32064 6092 32128
rect 6156 32064 6172 32128
rect 6236 32064 6252 32128
rect 6316 32064 6332 32128
rect 6396 32064 6404 32128
rect 6084 31040 6404 32064
rect 6084 30976 6092 31040
rect 6156 30976 6172 31040
rect 6236 30976 6252 31040
rect 6316 30976 6332 31040
rect 6396 30976 6404 31040
rect 6084 29952 6404 30976
rect 6084 29888 6092 29952
rect 6156 29888 6172 29952
rect 6236 29888 6252 29952
rect 6316 29888 6332 29952
rect 6396 29888 6404 29952
rect 6084 28864 6404 29888
rect 6084 28800 6092 28864
rect 6156 28800 6172 28864
rect 6236 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6404 28864
rect 6084 27776 6404 28800
rect 6084 27712 6092 27776
rect 6156 27712 6172 27776
rect 6236 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6404 27776
rect 6084 26688 6404 27712
rect 6084 26624 6092 26688
rect 6156 26624 6172 26688
rect 6236 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6404 26688
rect 6084 25600 6404 26624
rect 6084 25536 6092 25600
rect 6156 25536 6172 25600
rect 6236 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6404 25600
rect 6084 24512 6404 25536
rect 6499 25260 6565 25261
rect 6499 25196 6500 25260
rect 6564 25196 6565 25260
rect 6499 25195 6565 25196
rect 6084 24448 6092 24512
rect 6156 24448 6172 24512
rect 6236 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6404 24512
rect 6084 23424 6404 24448
rect 6084 23360 6092 23424
rect 6156 23360 6172 23424
rect 6236 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6404 23424
rect 6084 22336 6404 23360
rect 6084 22272 6092 22336
rect 6156 22272 6172 22336
rect 6236 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6404 22336
rect 6084 21248 6404 22272
rect 6084 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6404 21248
rect 6084 20160 6404 21184
rect 6084 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6404 20160
rect 6084 19072 6404 20096
rect 6084 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6404 19072
rect 6084 17984 6404 19008
rect 6084 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6404 17984
rect 6084 16896 6404 17920
rect 6502 17645 6562 25195
rect 6499 17644 6565 17645
rect 6499 17580 6500 17644
rect 6564 17580 6565 17644
rect 6499 17579 6565 17580
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6686 3501 6746 42603
rect 7797 42464 8117 43488
rect 7797 42400 7805 42464
rect 7869 42400 7885 42464
rect 7949 42400 7965 42464
rect 8029 42400 8045 42464
rect 8109 42400 8117 42464
rect 7419 41580 7485 41581
rect 7419 41516 7420 41580
rect 7484 41516 7485 41580
rect 7419 41515 7485 41516
rect 7235 31924 7301 31925
rect 7235 31860 7236 31924
rect 7300 31860 7301 31924
rect 7235 31859 7301 31860
rect 7238 23221 7298 31859
rect 7422 24037 7482 41515
rect 7797 41376 8117 42400
rect 7797 41312 7805 41376
rect 7869 41312 7885 41376
rect 7949 41312 7965 41376
rect 8029 41312 8045 41376
rect 8109 41312 8117 41376
rect 7797 40288 8117 41312
rect 7797 40224 7805 40288
rect 7869 40224 7885 40288
rect 7949 40224 7965 40288
rect 8029 40224 8045 40288
rect 8109 40224 8117 40288
rect 7797 39200 8117 40224
rect 9511 43008 9831 43568
rect 9511 42944 9519 43008
rect 9583 42944 9599 43008
rect 9663 42944 9679 43008
rect 9743 42944 9759 43008
rect 9823 42944 9831 43008
rect 9511 41920 9831 42944
rect 9511 41856 9519 41920
rect 9583 41856 9599 41920
rect 9663 41856 9679 41920
rect 9743 41856 9759 41920
rect 9823 41856 9831 41920
rect 9511 40832 9831 41856
rect 11224 43552 11544 43568
rect 11224 43488 11232 43552
rect 11296 43488 11312 43552
rect 11376 43488 11392 43552
rect 11456 43488 11472 43552
rect 11536 43488 11544 43552
rect 11224 42464 11544 43488
rect 11224 42400 11232 42464
rect 11296 42400 11312 42464
rect 11376 42400 11392 42464
rect 11456 42400 11472 42464
rect 11536 42400 11544 42464
rect 10915 41444 10981 41445
rect 10915 41380 10916 41444
rect 10980 41380 10981 41444
rect 10915 41379 10981 41380
rect 9511 40768 9519 40832
rect 9583 40768 9599 40832
rect 9663 40768 9679 40832
rect 9743 40768 9759 40832
rect 9823 40768 9831 40832
rect 9259 40084 9325 40085
rect 9259 40020 9260 40084
rect 9324 40020 9325 40084
rect 9259 40019 9325 40020
rect 7797 39136 7805 39200
rect 7869 39136 7885 39200
rect 7949 39136 7965 39200
rect 8029 39136 8045 39200
rect 8109 39136 8117 39200
rect 7797 38112 8117 39136
rect 7797 38048 7805 38112
rect 7869 38048 7885 38112
rect 7949 38048 7965 38112
rect 8029 38048 8045 38112
rect 8109 38048 8117 38112
rect 7797 37024 8117 38048
rect 7797 36960 7805 37024
rect 7869 36960 7885 37024
rect 7949 36960 7965 37024
rect 8029 36960 8045 37024
rect 8109 36960 8117 37024
rect 7797 35936 8117 36960
rect 7797 35872 7805 35936
rect 7869 35872 7885 35936
rect 7949 35872 7965 35936
rect 8029 35872 8045 35936
rect 8109 35872 8117 35936
rect 7797 34848 8117 35872
rect 7797 34784 7805 34848
rect 7869 34784 7885 34848
rect 7949 34784 7965 34848
rect 8029 34784 8045 34848
rect 8109 34784 8117 34848
rect 7797 33760 8117 34784
rect 7797 33696 7805 33760
rect 7869 33696 7885 33760
rect 7949 33696 7965 33760
rect 8029 33696 8045 33760
rect 8109 33696 8117 33760
rect 7797 32672 8117 33696
rect 8891 33284 8957 33285
rect 8891 33220 8892 33284
rect 8956 33220 8957 33284
rect 8891 33219 8957 33220
rect 7797 32608 7805 32672
rect 7869 32608 7885 32672
rect 7949 32608 7965 32672
rect 8029 32608 8045 32672
rect 8109 32608 8117 32672
rect 7797 31584 8117 32608
rect 7797 31520 7805 31584
rect 7869 31520 7885 31584
rect 7949 31520 7965 31584
rect 8029 31520 8045 31584
rect 8109 31520 8117 31584
rect 7797 30496 8117 31520
rect 7797 30432 7805 30496
rect 7869 30432 7885 30496
rect 7949 30432 7965 30496
rect 8029 30432 8045 30496
rect 8109 30432 8117 30496
rect 7797 29408 8117 30432
rect 7797 29344 7805 29408
rect 7869 29344 7885 29408
rect 7949 29344 7965 29408
rect 8029 29344 8045 29408
rect 8109 29344 8117 29408
rect 7797 28320 8117 29344
rect 7797 28256 7805 28320
rect 7869 28256 7885 28320
rect 7949 28256 7965 28320
rect 8029 28256 8045 28320
rect 8109 28256 8117 28320
rect 7797 27232 8117 28256
rect 7797 27168 7805 27232
rect 7869 27168 7885 27232
rect 7949 27168 7965 27232
rect 8029 27168 8045 27232
rect 8109 27168 8117 27232
rect 7797 26144 8117 27168
rect 7797 26080 7805 26144
rect 7869 26080 7885 26144
rect 7949 26080 7965 26144
rect 8029 26080 8045 26144
rect 8109 26080 8117 26144
rect 7797 25056 8117 26080
rect 7797 24992 7805 25056
rect 7869 24992 7885 25056
rect 7949 24992 7965 25056
rect 8029 24992 8045 25056
rect 8109 24992 8117 25056
rect 7419 24036 7485 24037
rect 7419 23972 7420 24036
rect 7484 23972 7485 24036
rect 7419 23971 7485 23972
rect 7797 23968 8117 24992
rect 7797 23904 7805 23968
rect 7869 23904 7885 23968
rect 7949 23904 7965 23968
rect 8029 23904 8045 23968
rect 8109 23904 8117 23968
rect 7419 23900 7485 23901
rect 7419 23836 7420 23900
rect 7484 23836 7485 23900
rect 7419 23835 7485 23836
rect 7235 23220 7301 23221
rect 7235 23156 7236 23220
rect 7300 23156 7301 23220
rect 7235 23155 7301 23156
rect 7422 18869 7482 23835
rect 7797 22880 8117 23904
rect 8894 23085 8954 33219
rect 9075 30836 9141 30837
rect 9075 30772 9076 30836
rect 9140 30772 9141 30836
rect 9075 30771 9141 30772
rect 8891 23084 8957 23085
rect 8891 23020 8892 23084
rect 8956 23020 8957 23084
rect 8891 23019 8957 23020
rect 7797 22816 7805 22880
rect 7869 22816 7885 22880
rect 7949 22816 7965 22880
rect 8029 22816 8045 22880
rect 8109 22816 8117 22880
rect 7603 21996 7669 21997
rect 7603 21932 7604 21996
rect 7668 21932 7669 21996
rect 7603 21931 7669 21932
rect 7419 18868 7485 18869
rect 7419 18804 7420 18868
rect 7484 18804 7485 18868
rect 7419 18803 7485 18804
rect 7419 18732 7485 18733
rect 7419 18668 7420 18732
rect 7484 18668 7485 18732
rect 7419 18667 7485 18668
rect 7422 12885 7482 18667
rect 7606 16557 7666 21931
rect 7797 21792 8117 22816
rect 8891 22540 8957 22541
rect 8891 22476 8892 22540
rect 8956 22476 8957 22540
rect 8891 22475 8957 22476
rect 7797 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8117 21792
rect 7797 20704 8117 21728
rect 7797 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8117 20704
rect 7797 19616 8117 20640
rect 7797 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8117 19616
rect 7797 18528 8117 19552
rect 7797 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8117 18528
rect 7797 17440 8117 18464
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7603 16556 7669 16557
rect 7603 16492 7604 16556
rect 7668 16492 7669 16556
rect 7603 16491 7669 16492
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 8894 15197 8954 22475
rect 9078 19549 9138 30771
rect 9262 22677 9322 40019
rect 9511 39744 9831 40768
rect 9511 39680 9519 39744
rect 9583 39680 9599 39744
rect 9663 39680 9679 39744
rect 9743 39680 9759 39744
rect 9823 39680 9831 39744
rect 9511 38656 9831 39680
rect 9511 38592 9519 38656
rect 9583 38592 9599 38656
rect 9663 38592 9679 38656
rect 9743 38592 9759 38656
rect 9823 38592 9831 38656
rect 9511 37568 9831 38592
rect 9511 37504 9519 37568
rect 9583 37504 9599 37568
rect 9663 37504 9679 37568
rect 9743 37504 9759 37568
rect 9823 37504 9831 37568
rect 9511 36480 9831 37504
rect 9511 36416 9519 36480
rect 9583 36416 9599 36480
rect 9663 36416 9679 36480
rect 9743 36416 9759 36480
rect 9823 36416 9831 36480
rect 9511 35392 9831 36416
rect 10547 36004 10613 36005
rect 10547 35940 10548 36004
rect 10612 35940 10613 36004
rect 10547 35939 10613 35940
rect 9511 35328 9519 35392
rect 9583 35328 9599 35392
rect 9663 35328 9679 35392
rect 9743 35328 9759 35392
rect 9823 35328 9831 35392
rect 9511 34304 9831 35328
rect 9511 34240 9519 34304
rect 9583 34240 9599 34304
rect 9663 34240 9679 34304
rect 9743 34240 9759 34304
rect 9823 34240 9831 34304
rect 9511 33216 9831 34240
rect 9511 33152 9519 33216
rect 9583 33152 9599 33216
rect 9663 33152 9679 33216
rect 9743 33152 9759 33216
rect 9823 33152 9831 33216
rect 9511 32128 9831 33152
rect 9511 32064 9519 32128
rect 9583 32064 9599 32128
rect 9663 32064 9679 32128
rect 9743 32064 9759 32128
rect 9823 32064 9831 32128
rect 9511 31040 9831 32064
rect 9511 30976 9519 31040
rect 9583 30976 9599 31040
rect 9663 30976 9679 31040
rect 9743 30976 9759 31040
rect 9823 30976 9831 31040
rect 9511 29952 9831 30976
rect 9511 29888 9519 29952
rect 9583 29888 9599 29952
rect 9663 29888 9679 29952
rect 9743 29888 9759 29952
rect 9823 29888 9831 29952
rect 9511 28864 9831 29888
rect 9511 28800 9519 28864
rect 9583 28800 9599 28864
rect 9663 28800 9679 28864
rect 9743 28800 9759 28864
rect 9823 28800 9831 28864
rect 9511 27776 9831 28800
rect 9511 27712 9519 27776
rect 9583 27712 9599 27776
rect 9663 27712 9679 27776
rect 9743 27712 9759 27776
rect 9823 27712 9831 27776
rect 9511 26688 9831 27712
rect 9511 26624 9519 26688
rect 9583 26624 9599 26688
rect 9663 26624 9679 26688
rect 9743 26624 9759 26688
rect 9823 26624 9831 26688
rect 9511 25600 9831 26624
rect 9511 25536 9519 25600
rect 9583 25536 9599 25600
rect 9663 25536 9679 25600
rect 9743 25536 9759 25600
rect 9823 25536 9831 25600
rect 9511 24512 9831 25536
rect 10550 25125 10610 35939
rect 10731 30700 10797 30701
rect 10731 30636 10732 30700
rect 10796 30636 10797 30700
rect 10731 30635 10797 30636
rect 10734 29613 10794 30635
rect 10731 29612 10797 29613
rect 10731 29548 10732 29612
rect 10796 29548 10797 29612
rect 10731 29547 10797 29548
rect 10547 25124 10613 25125
rect 10547 25060 10548 25124
rect 10612 25060 10613 25124
rect 10547 25059 10613 25060
rect 10547 24716 10613 24717
rect 10547 24652 10548 24716
rect 10612 24652 10613 24716
rect 10547 24651 10613 24652
rect 9511 24448 9519 24512
rect 9583 24448 9599 24512
rect 9663 24448 9679 24512
rect 9743 24448 9759 24512
rect 9823 24448 9831 24512
rect 9511 23424 9831 24448
rect 9511 23360 9519 23424
rect 9583 23360 9599 23424
rect 9663 23360 9679 23424
rect 9743 23360 9759 23424
rect 9823 23360 9831 23424
rect 9259 22676 9325 22677
rect 9259 22612 9260 22676
rect 9324 22612 9325 22676
rect 9259 22611 9325 22612
rect 9075 19548 9141 19549
rect 9075 19484 9076 19548
rect 9140 19484 9141 19548
rect 9075 19483 9141 19484
rect 9262 16557 9322 22611
rect 9511 22336 9831 23360
rect 9511 22272 9519 22336
rect 9583 22272 9599 22336
rect 9663 22272 9679 22336
rect 9743 22272 9759 22336
rect 9823 22272 9831 22336
rect 9511 21248 9831 22272
rect 9995 21724 10061 21725
rect 9995 21660 9996 21724
rect 10060 21660 10061 21724
rect 9995 21659 10061 21660
rect 9511 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9831 21248
rect 9511 20160 9831 21184
rect 9511 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9831 20160
rect 9511 19072 9831 20096
rect 9998 19549 10058 21659
rect 9995 19548 10061 19549
rect 9995 19484 9996 19548
rect 10060 19484 10061 19548
rect 9995 19483 10061 19484
rect 9511 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9831 19072
rect 9511 17984 9831 19008
rect 9511 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9831 17984
rect 9511 16896 9831 17920
rect 10550 17781 10610 24651
rect 10734 18733 10794 29547
rect 10731 18732 10797 18733
rect 10731 18668 10732 18732
rect 10796 18668 10797 18732
rect 10731 18667 10797 18668
rect 10547 17780 10613 17781
rect 10547 17716 10548 17780
rect 10612 17716 10613 17780
rect 10547 17715 10613 17716
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 9259 16556 9325 16557
rect 9259 16492 9260 16556
rect 9324 16492 9325 16556
rect 9259 16491 9325 16492
rect 9511 15808 9831 16832
rect 10547 16420 10613 16421
rect 10547 16356 10548 16420
rect 10612 16356 10613 16420
rect 10547 16355 10613 16356
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 8891 15196 8957 15197
rect 8891 15132 8892 15196
rect 8956 15132 8957 15196
rect 8891 15131 8957 15132
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7419 12884 7485 12885
rect 7419 12820 7420 12884
rect 7484 12820 7485 12884
rect 7419 12819 7485 12820
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 6683 3500 6749 3501
rect 6683 3436 6684 3500
rect 6748 3436 6749 3500
rect 6683 3435 6749 3436
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 1664 6404 2688
rect 6084 1600 6092 1664
rect 6156 1600 6172 1664
rect 6236 1600 6252 1664
rect 6316 1600 6332 1664
rect 6396 1600 6404 1664
rect 4843 1324 4909 1325
rect 4843 1260 4844 1324
rect 4908 1260 4909 1324
rect 4843 1259 4909 1260
rect 5395 1324 5461 1325
rect 5395 1260 5396 1324
rect 5460 1260 5461 1324
rect 5395 1259 5461 1260
rect 4370 1056 4378 1120
rect 4442 1056 4458 1120
rect 4522 1056 4538 1120
rect 4602 1056 4618 1120
rect 4682 1056 4690 1120
rect 4370 1040 4690 1056
rect 6084 1040 6404 1600
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 1120 8117 2144
rect 7797 1056 7805 1120
rect 7869 1056 7885 1120
rect 7949 1056 7965 1120
rect 8029 1056 8045 1120
rect 8109 1056 8117 1120
rect 7797 1040 8117 1056
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 9511 13632 9831 14656
rect 10550 13837 10610 16355
rect 10734 14381 10794 18667
rect 10731 14380 10797 14381
rect 10731 14316 10732 14380
rect 10796 14316 10797 14380
rect 10731 14315 10797 14316
rect 10547 13836 10613 13837
rect 10547 13772 10548 13836
rect 10612 13772 10613 13836
rect 10547 13771 10613 13772
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 1664 9831 2688
rect 10918 2685 10978 41379
rect 11224 41376 11544 42400
rect 11224 41312 11232 41376
rect 11296 41312 11312 41376
rect 11376 41312 11392 41376
rect 11456 41312 11472 41376
rect 11536 41312 11544 41376
rect 11224 40288 11544 41312
rect 11224 40224 11232 40288
rect 11296 40224 11312 40288
rect 11376 40224 11392 40288
rect 11456 40224 11472 40288
rect 11536 40224 11544 40288
rect 11224 39200 11544 40224
rect 11224 39136 11232 39200
rect 11296 39136 11312 39200
rect 11376 39136 11392 39200
rect 11456 39136 11472 39200
rect 11536 39136 11544 39200
rect 11224 38112 11544 39136
rect 11224 38048 11232 38112
rect 11296 38048 11312 38112
rect 11376 38048 11392 38112
rect 11456 38048 11472 38112
rect 11536 38048 11544 38112
rect 11224 37024 11544 38048
rect 11224 36960 11232 37024
rect 11296 36960 11312 37024
rect 11376 36960 11392 37024
rect 11456 36960 11472 37024
rect 11536 36960 11544 37024
rect 11224 35936 11544 36960
rect 11224 35872 11232 35936
rect 11296 35872 11312 35936
rect 11376 35872 11392 35936
rect 11456 35872 11472 35936
rect 11536 35872 11544 35936
rect 11224 34848 11544 35872
rect 11224 34784 11232 34848
rect 11296 34784 11312 34848
rect 11376 34784 11392 34848
rect 11456 34784 11472 34848
rect 11536 34784 11544 34848
rect 11224 33760 11544 34784
rect 12938 43008 13258 43568
rect 12938 42944 12946 43008
rect 13010 42944 13026 43008
rect 13090 42944 13106 43008
rect 13170 42944 13186 43008
rect 13250 42944 13258 43008
rect 12938 41920 13258 42944
rect 12938 41856 12946 41920
rect 13010 41856 13026 41920
rect 13090 41856 13106 41920
rect 13170 41856 13186 41920
rect 13250 41856 13258 41920
rect 12938 40832 13258 41856
rect 12938 40768 12946 40832
rect 13010 40768 13026 40832
rect 13090 40768 13106 40832
rect 13170 40768 13186 40832
rect 13250 40768 13258 40832
rect 12938 39744 13258 40768
rect 12938 39680 12946 39744
rect 13010 39680 13026 39744
rect 13090 39680 13106 39744
rect 13170 39680 13186 39744
rect 13250 39680 13258 39744
rect 12938 38656 13258 39680
rect 12938 38592 12946 38656
rect 13010 38592 13026 38656
rect 13090 38592 13106 38656
rect 13170 38592 13186 38656
rect 13250 38592 13258 38656
rect 12938 37568 13258 38592
rect 12938 37504 12946 37568
rect 13010 37504 13026 37568
rect 13090 37504 13106 37568
rect 13170 37504 13186 37568
rect 13250 37504 13258 37568
rect 12938 36480 13258 37504
rect 12938 36416 12946 36480
rect 13010 36416 13026 36480
rect 13090 36416 13106 36480
rect 13170 36416 13186 36480
rect 13250 36416 13258 36480
rect 12938 35392 13258 36416
rect 12938 35328 12946 35392
rect 13010 35328 13026 35392
rect 13090 35328 13106 35392
rect 13170 35328 13186 35392
rect 13250 35328 13258 35392
rect 12938 34304 13258 35328
rect 12938 34240 12946 34304
rect 13010 34240 13026 34304
rect 13090 34240 13106 34304
rect 13170 34240 13186 34304
rect 13250 34240 13258 34304
rect 11651 33964 11717 33965
rect 11651 33900 11652 33964
rect 11716 33900 11717 33964
rect 11651 33899 11717 33900
rect 11224 33696 11232 33760
rect 11296 33696 11312 33760
rect 11376 33696 11392 33760
rect 11456 33696 11472 33760
rect 11536 33696 11544 33760
rect 11224 32672 11544 33696
rect 11224 32608 11232 32672
rect 11296 32608 11312 32672
rect 11376 32608 11392 32672
rect 11456 32608 11472 32672
rect 11536 32608 11544 32672
rect 11224 31584 11544 32608
rect 11224 31520 11232 31584
rect 11296 31520 11312 31584
rect 11376 31520 11392 31584
rect 11456 31520 11472 31584
rect 11536 31520 11544 31584
rect 11224 30496 11544 31520
rect 11224 30432 11232 30496
rect 11296 30432 11312 30496
rect 11376 30432 11392 30496
rect 11456 30432 11472 30496
rect 11536 30432 11544 30496
rect 11224 29408 11544 30432
rect 11224 29344 11232 29408
rect 11296 29344 11312 29408
rect 11376 29344 11392 29408
rect 11456 29344 11472 29408
rect 11536 29344 11544 29408
rect 11224 28320 11544 29344
rect 11654 29069 11714 33899
rect 12938 33216 13258 34240
rect 14651 43552 14971 43568
rect 14651 43488 14659 43552
rect 14723 43488 14739 43552
rect 14803 43488 14819 43552
rect 14883 43488 14899 43552
rect 14963 43488 14971 43552
rect 14651 42464 14971 43488
rect 14651 42400 14659 42464
rect 14723 42400 14739 42464
rect 14803 42400 14819 42464
rect 14883 42400 14899 42464
rect 14963 42400 14971 42464
rect 14651 41376 14971 42400
rect 14651 41312 14659 41376
rect 14723 41312 14739 41376
rect 14803 41312 14819 41376
rect 14883 41312 14899 41376
rect 14963 41312 14971 41376
rect 14651 40288 14971 41312
rect 14651 40224 14659 40288
rect 14723 40224 14739 40288
rect 14803 40224 14819 40288
rect 14883 40224 14899 40288
rect 14963 40224 14971 40288
rect 14651 39200 14971 40224
rect 14651 39136 14659 39200
rect 14723 39136 14739 39200
rect 14803 39136 14819 39200
rect 14883 39136 14899 39200
rect 14963 39136 14971 39200
rect 14651 38112 14971 39136
rect 14651 38048 14659 38112
rect 14723 38048 14739 38112
rect 14803 38048 14819 38112
rect 14883 38048 14899 38112
rect 14963 38048 14971 38112
rect 14651 37024 14971 38048
rect 14651 36960 14659 37024
rect 14723 36960 14739 37024
rect 14803 36960 14819 37024
rect 14883 36960 14899 37024
rect 14963 36960 14971 37024
rect 14651 35936 14971 36960
rect 14651 35872 14659 35936
rect 14723 35872 14739 35936
rect 14803 35872 14819 35936
rect 14883 35872 14899 35936
rect 14963 35872 14971 35936
rect 14651 34848 14971 35872
rect 14651 34784 14659 34848
rect 14723 34784 14739 34848
rect 14803 34784 14819 34848
rect 14883 34784 14899 34848
rect 14963 34784 14971 34848
rect 14651 33760 14971 34784
rect 14651 33696 14659 33760
rect 14723 33696 14739 33760
rect 14803 33696 14819 33760
rect 14883 33696 14899 33760
rect 14963 33696 14971 33760
rect 13491 33692 13557 33693
rect 13491 33628 13492 33692
rect 13556 33628 13557 33692
rect 13491 33627 13557 33628
rect 12938 33152 12946 33216
rect 13010 33152 13026 33216
rect 13090 33152 13106 33216
rect 13170 33152 13186 33216
rect 13250 33152 13258 33216
rect 12755 32740 12821 32741
rect 12755 32676 12756 32740
rect 12820 32676 12821 32740
rect 12755 32675 12821 32676
rect 12571 32604 12637 32605
rect 12571 32540 12572 32604
rect 12636 32540 12637 32604
rect 12571 32539 12637 32540
rect 12574 30157 12634 32539
rect 12571 30156 12637 30157
rect 12571 30092 12572 30156
rect 12636 30092 12637 30156
rect 12571 30091 12637 30092
rect 11651 29068 11717 29069
rect 11651 29004 11652 29068
rect 11716 29004 11717 29068
rect 11651 29003 11717 29004
rect 11224 28256 11232 28320
rect 11296 28256 11312 28320
rect 11376 28256 11392 28320
rect 11456 28256 11472 28320
rect 11536 28256 11544 28320
rect 11224 27232 11544 28256
rect 11224 27168 11232 27232
rect 11296 27168 11312 27232
rect 11376 27168 11392 27232
rect 11456 27168 11472 27232
rect 11536 27168 11544 27232
rect 11224 26144 11544 27168
rect 11224 26080 11232 26144
rect 11296 26080 11312 26144
rect 11376 26080 11392 26144
rect 11456 26080 11472 26144
rect 11536 26080 11544 26144
rect 11224 25056 11544 26080
rect 11224 24992 11232 25056
rect 11296 24992 11312 25056
rect 11376 24992 11392 25056
rect 11456 24992 11472 25056
rect 11536 24992 11544 25056
rect 11224 23968 11544 24992
rect 11224 23904 11232 23968
rect 11296 23904 11312 23968
rect 11376 23904 11392 23968
rect 11456 23904 11472 23968
rect 11536 23904 11544 23968
rect 11224 22880 11544 23904
rect 12574 23085 12634 30091
rect 12758 29885 12818 32675
rect 12938 32128 13258 33152
rect 12938 32064 12946 32128
rect 13010 32064 13026 32128
rect 13090 32064 13106 32128
rect 13170 32064 13186 32128
rect 13250 32064 13258 32128
rect 12938 31040 13258 32064
rect 12938 30976 12946 31040
rect 13010 30976 13026 31040
rect 13090 30976 13106 31040
rect 13170 30976 13186 31040
rect 13250 30976 13258 31040
rect 12938 29952 13258 30976
rect 12938 29888 12946 29952
rect 13010 29888 13026 29952
rect 13090 29888 13106 29952
rect 13170 29888 13186 29952
rect 13250 29888 13258 29952
rect 12755 29884 12821 29885
rect 12755 29820 12756 29884
rect 12820 29820 12821 29884
rect 12755 29819 12821 29820
rect 12938 28864 13258 29888
rect 13494 29205 13554 33627
rect 14651 32672 14971 33696
rect 14651 32608 14659 32672
rect 14723 32608 14739 32672
rect 14803 32608 14819 32672
rect 14883 32608 14899 32672
rect 14963 32608 14971 32672
rect 14043 31788 14109 31789
rect 14043 31724 14044 31788
rect 14108 31724 14109 31788
rect 14043 31723 14109 31724
rect 13491 29204 13557 29205
rect 13491 29140 13492 29204
rect 13556 29140 13557 29204
rect 13491 29139 13557 29140
rect 12938 28800 12946 28864
rect 13010 28800 13026 28864
rect 13090 28800 13106 28864
rect 13170 28800 13186 28864
rect 13250 28800 13258 28864
rect 12755 28796 12821 28797
rect 12755 28732 12756 28796
rect 12820 28732 12821 28796
rect 12755 28731 12821 28732
rect 12758 28525 12818 28731
rect 12755 28524 12821 28525
rect 12755 28460 12756 28524
rect 12820 28460 12821 28524
rect 12755 28459 12821 28460
rect 12938 27776 13258 28800
rect 12938 27712 12946 27776
rect 13010 27712 13026 27776
rect 13090 27712 13106 27776
rect 13170 27712 13186 27776
rect 13250 27712 13258 27776
rect 12938 26688 13258 27712
rect 12938 26624 12946 26688
rect 13010 26624 13026 26688
rect 13090 26624 13106 26688
rect 13170 26624 13186 26688
rect 13250 26624 13258 26688
rect 12938 25600 13258 26624
rect 12938 25536 12946 25600
rect 13010 25536 13026 25600
rect 13090 25536 13106 25600
rect 13170 25536 13186 25600
rect 13250 25536 13258 25600
rect 12938 24512 13258 25536
rect 13494 24717 13554 29139
rect 13859 28252 13925 28253
rect 13859 28188 13860 28252
rect 13924 28188 13925 28252
rect 13859 28187 13925 28188
rect 13675 27436 13741 27437
rect 13675 27372 13676 27436
rect 13740 27372 13741 27436
rect 13675 27371 13741 27372
rect 13491 24716 13557 24717
rect 13491 24652 13492 24716
rect 13556 24652 13557 24716
rect 13491 24651 13557 24652
rect 12938 24448 12946 24512
rect 13010 24448 13026 24512
rect 13090 24448 13106 24512
rect 13170 24448 13186 24512
rect 13250 24448 13258 24512
rect 12938 23424 13258 24448
rect 12938 23360 12946 23424
rect 13010 23360 13026 23424
rect 13090 23360 13106 23424
rect 13170 23360 13186 23424
rect 13250 23360 13258 23424
rect 11651 23084 11717 23085
rect 11651 23020 11652 23084
rect 11716 23020 11717 23084
rect 11651 23019 11717 23020
rect 12571 23084 12637 23085
rect 12571 23020 12572 23084
rect 12636 23020 12637 23084
rect 12571 23019 12637 23020
rect 11224 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11392 22880
rect 11456 22816 11472 22880
rect 11536 22816 11544 22880
rect 11224 21792 11544 22816
rect 11224 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11544 21792
rect 11224 20704 11544 21728
rect 11224 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11544 20704
rect 11224 19616 11544 20640
rect 11224 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11544 19616
rect 11224 18528 11544 19552
rect 11224 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11544 18528
rect 11224 17440 11544 18464
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11654 17101 11714 23019
rect 11835 22676 11901 22677
rect 11835 22612 11836 22676
rect 11900 22612 11901 22676
rect 11835 22611 11901 22612
rect 11838 19005 11898 22611
rect 12203 21180 12269 21181
rect 12203 21116 12204 21180
rect 12268 21116 12269 21180
rect 12203 21115 12269 21116
rect 11835 19004 11901 19005
rect 11835 18940 11836 19004
rect 11900 18940 11901 19004
rect 11835 18939 11901 18940
rect 11835 17644 11901 17645
rect 11835 17580 11836 17644
rect 11900 17580 11901 17644
rect 11835 17579 11901 17580
rect 11651 17100 11717 17101
rect 11651 17036 11652 17100
rect 11716 17036 11717 17100
rect 11651 17035 11717 17036
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 11224 8736 11544 9760
rect 11651 9756 11717 9757
rect 11651 9692 11652 9756
rect 11716 9692 11717 9756
rect 11651 9691 11717 9692
rect 11654 9349 11714 9691
rect 11651 9348 11717 9349
rect 11651 9284 11652 9348
rect 11716 9284 11717 9348
rect 11651 9283 11717 9284
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 10915 2684 10981 2685
rect 10915 2620 10916 2684
rect 10980 2620 10981 2684
rect 10915 2619 10981 2620
rect 9511 1600 9519 1664
rect 9583 1600 9599 1664
rect 9663 1600 9679 1664
rect 9743 1600 9759 1664
rect 9823 1600 9831 1664
rect 9511 1040 9831 1600
rect 11224 2208 11544 3232
rect 11838 2685 11898 17579
rect 12206 16829 12266 21115
rect 12574 18869 12634 23019
rect 12938 22336 13258 23360
rect 12938 22272 12946 22336
rect 13010 22272 13026 22336
rect 13090 22272 13106 22336
rect 13170 22272 13186 22336
rect 13250 22272 13258 22336
rect 12755 22132 12821 22133
rect 12755 22068 12756 22132
rect 12820 22068 12821 22132
rect 12755 22067 12821 22068
rect 12571 18868 12637 18869
rect 12571 18804 12572 18868
rect 12636 18804 12637 18868
rect 12571 18803 12637 18804
rect 12203 16828 12269 16829
rect 12203 16764 12204 16828
rect 12268 16764 12269 16828
rect 12203 16763 12269 16764
rect 12758 15333 12818 22067
rect 12938 21248 13258 22272
rect 12938 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13258 21248
rect 12938 20160 13258 21184
rect 12938 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13258 20160
rect 12938 19072 13258 20096
rect 13678 19957 13738 27371
rect 13675 19956 13741 19957
rect 13675 19892 13676 19956
rect 13740 19892 13741 19956
rect 13675 19891 13741 19892
rect 12938 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13258 19072
rect 12938 17984 13258 19008
rect 12938 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13258 17984
rect 12938 16896 13258 17920
rect 13862 17917 13922 28187
rect 13859 17916 13925 17917
rect 13859 17852 13860 17916
rect 13924 17852 13925 17916
rect 13859 17851 13925 17852
rect 13491 17372 13557 17373
rect 13491 17308 13492 17372
rect 13556 17308 13557 17372
rect 13491 17307 13557 17308
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12938 15808 13258 16832
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 12755 15332 12821 15333
rect 12755 15268 12756 15332
rect 12820 15268 12821 15332
rect 12755 15267 12821 15268
rect 12755 15196 12821 15197
rect 12755 15132 12756 15196
rect 12820 15132 12821 15196
rect 12755 15131 12821 15132
rect 12758 10029 12818 15131
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 13494 11797 13554 17307
rect 14046 16693 14106 31723
rect 14651 31584 14971 32608
rect 14651 31520 14659 31584
rect 14723 31520 14739 31584
rect 14803 31520 14819 31584
rect 14883 31520 14899 31584
rect 14963 31520 14971 31584
rect 14651 30496 14971 31520
rect 14651 30432 14659 30496
rect 14723 30432 14739 30496
rect 14803 30432 14819 30496
rect 14883 30432 14899 30496
rect 14963 30432 14971 30496
rect 14651 29408 14971 30432
rect 14651 29344 14659 29408
rect 14723 29344 14739 29408
rect 14803 29344 14819 29408
rect 14883 29344 14899 29408
rect 14963 29344 14971 29408
rect 14651 28320 14971 29344
rect 14651 28256 14659 28320
rect 14723 28256 14739 28320
rect 14803 28256 14819 28320
rect 14883 28256 14899 28320
rect 14963 28256 14971 28320
rect 14651 27232 14971 28256
rect 14651 27168 14659 27232
rect 14723 27168 14739 27232
rect 14803 27168 14819 27232
rect 14883 27168 14899 27232
rect 14963 27168 14971 27232
rect 14651 26144 14971 27168
rect 14651 26080 14659 26144
rect 14723 26080 14739 26144
rect 14803 26080 14819 26144
rect 14883 26080 14899 26144
rect 14963 26080 14971 26144
rect 14651 25056 14971 26080
rect 14651 24992 14659 25056
rect 14723 24992 14739 25056
rect 14803 24992 14819 25056
rect 14883 24992 14899 25056
rect 14963 24992 14971 25056
rect 14651 23968 14971 24992
rect 14651 23904 14659 23968
rect 14723 23904 14739 23968
rect 14803 23904 14819 23968
rect 14883 23904 14899 23968
rect 14963 23904 14971 23968
rect 14651 22880 14971 23904
rect 14651 22816 14659 22880
rect 14723 22816 14739 22880
rect 14803 22816 14819 22880
rect 14883 22816 14899 22880
rect 14963 22816 14971 22880
rect 14651 21792 14971 22816
rect 14651 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14971 21792
rect 14651 20704 14971 21728
rect 14651 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14971 20704
rect 14651 19616 14971 20640
rect 14651 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14971 19616
rect 14651 18528 14971 19552
rect 14651 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14971 18528
rect 14227 17508 14293 17509
rect 14227 17444 14228 17508
rect 14292 17444 14293 17508
rect 14227 17443 14293 17444
rect 14043 16692 14109 16693
rect 14043 16628 14044 16692
rect 14108 16628 14109 16692
rect 14043 16627 14109 16628
rect 13675 14924 13741 14925
rect 13675 14860 13676 14924
rect 13740 14860 13741 14924
rect 13675 14859 13741 14860
rect 13678 11933 13738 14859
rect 14046 12205 14106 16627
rect 14230 13837 14290 17443
rect 14651 17440 14971 18464
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14227 13836 14293 13837
rect 14227 13772 14228 13836
rect 14292 13772 14293 13836
rect 14227 13771 14293 13772
rect 14651 13088 14971 14112
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14043 12204 14109 12205
rect 14043 12140 14044 12204
rect 14108 12140 14109 12204
rect 14043 12139 14109 12140
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 13675 11932 13741 11933
rect 13675 11868 13676 11932
rect 13740 11868 13741 11932
rect 13675 11867 13741 11868
rect 13491 11796 13557 11797
rect 13491 11732 13492 11796
rect 13556 11732 13557 11796
rect 13491 11731 13557 11732
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12755 10028 12821 10029
rect 12755 9964 12756 10028
rect 12820 9964 12821 10028
rect 12755 9963 12821 9964
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12203 9076 12269 9077
rect 12203 9012 12204 9076
rect 12268 9012 12269 9076
rect 12203 9011 12269 9012
rect 12206 8669 12266 9011
rect 12203 8668 12269 8669
rect 12203 8604 12204 8668
rect 12268 8604 12269 8668
rect 12203 8603 12269 8604
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 11835 2684 11901 2685
rect 11835 2620 11836 2684
rect 11900 2620 11901 2684
rect 11835 2619 11901 2620
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 1120 11544 2144
rect 11224 1056 11232 1120
rect 11296 1056 11312 1120
rect 11376 1056 11392 1120
rect 11456 1056 11472 1120
rect 11536 1056 11544 1120
rect 11224 1040 11544 1056
rect 12938 1664 13258 2688
rect 12938 1600 12946 1664
rect 13010 1600 13026 1664
rect 13090 1600 13106 1664
rect 13170 1600 13186 1664
rect 13250 1600 13258 1664
rect 12938 1040 13258 1600
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 1120 14971 2144
rect 14651 1056 14659 1120
rect 14723 1056 14739 1120
rect 14803 1056 14819 1120
rect 14883 1056 14899 1120
rect 14963 1056 14971 1120
rect 14651 1040 14971 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9844 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform -1 0 13800 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0__0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1__0_
timestamp 1688980957
transform 1 0 13524 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2__0_
timestamp 1688980957
transform 1 0 10672 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3__0_
timestamp 1688980957
transform 1 0 10948 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4__0_
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5__0_
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6__0_
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7__0_
timestamp 1688980957
transform 1 0 9936 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8__0_
timestamp 1688980957
transform 1 0 11224 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9__0_
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10__0_
timestamp 1688980957
transform 1 0 10396 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11__0_
timestamp 1688980957
transform 1 0 12052 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12__0_
timestamp 1688980957
transform 1 0 10488 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13__0_
timestamp 1688980957
transform 1 0 12328 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14__0_
timestamp 1688980957
transform 1 0 10212 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15__0_
timestamp 1688980957
transform 1 0 10948 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16__0_
timestamp 1688980957
transform 1 0 12604 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17__0_
timestamp 1688980957
transform 1 0 12052 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18__0_
timestamp 1688980957
transform 1 0 9292 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19__0_
timestamp 1688980957
transform 1 0 8372 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20__0_
timestamp 1688980957
transform 1 0 11776 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21__0_
timestamp 1688980957
transform 1 0 11500 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22__0_
timestamp 1688980957
transform 1 0 12880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23__0_
timestamp 1688980957
transform 1 0 11868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24__0_
timestamp 1688980957
transform 1 0 12328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25__0_
timestamp 1688980957
transform 1 0 13248 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26__0_
timestamp 1688980957
transform 1 0 10764 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27__0_
timestamp 1688980957
transform 1 0 11776 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28__0_
timestamp 1688980957
transform 1 0 12696 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29__0_
timestamp 1688980957
transform 1 0 12696 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30__0_
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31__0_
timestamp 1688980957
transform 1 0 9200 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0__0_
timestamp 1688980957
transform 1 0 10948 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1__0_
timestamp 1688980957
transform 1 0 10488 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2__0_
timestamp 1688980957
transform 1 0 10764 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3__0_
timestamp 1688980957
transform 1 0 11040 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4__0_
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5__0_
timestamp 1688980957
transform 1 0 11500 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6__0_
timestamp 1688980957
transform 1 0 9476 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7__0_
timestamp 1688980957
transform 1 0 10488 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8__0_
timestamp 1688980957
transform 1 0 11592 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9__0_
timestamp 1688980957
transform 1 0 10672 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10__0_
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11__0_
timestamp 1688980957
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12__0_
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13__0_
timestamp 1688980957
transform 1 0 12420 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14__0_
timestamp 1688980957
transform 1 0 11776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15__0_
timestamp 1688980957
transform 1 0 11224 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16__0_
timestamp 1688980957
transform 1 0 12696 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17__0_
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18__0_
timestamp 1688980957
transform 1 0 10120 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19__0_
timestamp 1688980957
transform 1 0 9108 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20__0_
timestamp 1688980957
transform 1 0 13156 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21__0_
timestamp 1688980957
transform 1 0 12144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22__0_
timestamp 1688980957
transform 1 0 12604 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23__0_
timestamp 1688980957
transform 1 0 12972 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24__0_
timestamp 1688980957
transform 1 0 12972 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25__0_
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26__0_
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27__0_
timestamp 1688980957
transform 1 0 12420 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28__0_
timestamp 1688980957
transform 1 0 12696 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29__0_
timestamp 1688980957
transform 1 0 12972 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30__0_
timestamp 1688980957
transform 1 0 9476 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31__0_
timestamp 1688980957
transform 1 0 10028 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3220 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_39
timestamp 1688980957
transform 1 0 4692 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_47
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_62
timestamp 1688980957
transform 1 0 6808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_66
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_70
timestamp 1688980957
transform 1 0 7544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_74
timestamp 1688980957
transform 1 0 7912 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_78 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_88 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_94
timestamp 1688980957
transform 1 0 9752 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_98
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_102
timestamp 1688980957
transform 1 0 10488 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_106
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_118
timestamp 1688980957
transform 1 0 11960 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_122
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 1688980957
transform 1 0 14444 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_31 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_43
timestamp 1688980957
transform 1 0 5060 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_53
timestamp 1688980957
transform 1 0 5980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_61
timestamp 1688980957
transform 1 0 6716 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_77
timestamp 1688980957
transform 1 0 8188 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_84
timestamp 1688980957
transform 1 0 8832 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_92
timestamp 1688980957
transform 1 0 9568 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_96
timestamp 1688980957
transform 1 0 9936 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_101
timestamp 1688980957
transform 1 0 10396 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 1688980957
transform 1 0 11132 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_117
timestamp 1688980957
transform 1 0 11868 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_132
timestamp 1688980957
transform 1 0 13248 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_145
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_133
timestamp 1688980957
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_129
timestamp 1688980957
transform 1 0 12972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_145
timestamp 1688980957
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_143
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1688980957
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_118
timestamp 1688980957
transform 1 0 11960 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_124
timestamp 1688980957
transform 1 0 12512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_145
timestamp 1688980957
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_21
timestamp 1688980957
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_45
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1688980957
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_75
timestamp 1688980957
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 1688980957
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_145
timestamp 1688980957
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_9
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_16
timestamp 1688980957
transform 1 0 2576 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_105
timestamp 1688980957
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_18
timestamp 1688980957
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_42
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_75
timestamp 1688980957
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_134
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_17
timestamp 1688980957
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1688980957
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1688980957
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1688980957
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_42
timestamp 1688980957
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1688980957
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1688980957
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_61
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_103
timestamp 1688980957
transform 1 0 10580 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_129
timestamp 1688980957
transform 1 0 12972 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_135
timestamp 1688980957
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_12
timestamp 1688980957
transform 1 0 2208 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_24
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_36
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_48
timestamp 1688980957
transform 1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_52
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_61
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_66
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_89
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_143
timestamp 1688980957
transform 1 0 14260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_18
timestamp 1688980957
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_130
timestamp 1688980957
transform 1 0 13064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_21
timestamp 1688980957
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_33
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_45
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_61
timestamp 1688980957
transform 1 0 6716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_73
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_82
timestamp 1688980957
transform 1 0 8648 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_90
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_134
timestamp 1688980957
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_9
timestamp 1688980957
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_16
timestamp 1688980957
transform 1 0 2576 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_64
timestamp 1688980957
transform 1 0 6992 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_76
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_8
timestamp 1688980957
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_20
timestamp 1688980957
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_32
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_44
timestamp 1688980957
transform 1 0 5152 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_83
timestamp 1688980957
transform 1 0 8740 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_95
timestamp 1688980957
transform 1 0 9844 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_107
timestamp 1688980957
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_126
timestamp 1688980957
transform 1 0 12696 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_145
timestamp 1688980957
transform 1 0 14444 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_9
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_21
timestamp 1688980957
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_101
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_105
timestamp 1688980957
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_21
timestamp 1688980957
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_33
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_66
timestamp 1688980957
transform 1 0 7176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_103
timestamp 1688980957
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_12
timestamp 1688980957
transform 1 0 2208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp 1688980957
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_74
timestamp 1688980957
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1688980957
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 1688980957
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_30
timestamp 1688980957
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_21
timestamp 1688980957
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_100
timestamp 1688980957
transform 1 0 10304 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_112
timestamp 1688980957
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_12
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_24
timestamp 1688980957
transform 1 0 3312 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_36
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_48
timestamp 1688980957
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_102
timestamp 1688980957
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1688980957
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_18
timestamp 1688980957
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1688980957
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_49
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_122
timestamp 1688980957
transform 1 0 12328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_12
timestamp 1688980957
transform 1 0 2208 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_24
timestamp 1688980957
transform 1 0 3312 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_36
timestamp 1688980957
transform 1 0 4416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_48
timestamp 1688980957
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_75
timestamp 1688980957
transform 1 0 8004 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_87
timestamp 1688980957
transform 1 0 9108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_119
timestamp 1688980957
transform 1 0 12052 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_144
timestamp 1688980957
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_10
timestamp 1688980957
transform 1 0 2024 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_22
timestamp 1688980957
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_62
timestamp 1688980957
transform 1 0 6808 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_74
timestamp 1688980957
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_18
timestamp 1688980957
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_30
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_42
timestamp 1688980957
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_65
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_102
timestamp 1688980957
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1688980957
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_18
timestamp 1688980957
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_76
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1688980957
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_7
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_19
timestamp 1688980957
transform 1 0 2852 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_31
timestamp 1688980957
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_43
timestamp 1688980957
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_86
timestamp 1688980957
transform 1 0 9016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_90
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_129
timestamp 1688980957
transform 1 0 12972 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_7
timestamp 1688980957
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_70
timestamp 1688980957
transform 1 0 7544 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_82
timestamp 1688980957
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_89
timestamp 1688980957
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_105
timestamp 1688980957
transform 1 0 10764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_145
timestamp 1688980957
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_7
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_19
timestamp 1688980957
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_31
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_61
timestamp 1688980957
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_77
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_96
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_108
timestamp 1688980957
transform 1 0 11040 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_117
timestamp 1688980957
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_124
timestamp 1688980957
transform 1 0 12512 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_66
timestamp 1688980957
transform 1 0 7176 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_73
timestamp 1688980957
transform 1 0 7820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_144
timestamp 1688980957
transform 1 0 14352 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_7
timestamp 1688980957
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_19
timestamp 1688980957
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_31
timestamp 1688980957
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_43
timestamp 1688980957
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_61
timestamp 1688980957
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_72
timestamp 1688980957
transform 1 0 7728 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_89
timestamp 1688980957
transform 1 0 9292 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_101
timestamp 1688980957
transform 1 0 10396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 1688980957
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_124
timestamp 1688980957
transform 1 0 12512 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_141
timestamp 1688980957
transform 1 0 14076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 1688980957
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_49
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_106
timestamp 1688980957
transform 1 0 10856 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_145
timestamp 1688980957
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_61
timestamp 1688980957
transform 1 0 6716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_70
timestamp 1688980957
transform 1 0 7544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_76
timestamp 1688980957
transform 1 0 8096 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_135
timestamp 1688980957
transform 1 0 13524 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_142
timestamp 1688980957
transform 1 0 14168 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_13
timestamp 1688980957
transform 1 0 2300 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_21
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_25
timestamp 1688980957
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_78
timestamp 1688980957
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_93
timestamp 1688980957
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_145
timestamp 1688980957
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_7
timestamp 1688980957
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_19
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_31
timestamp 1688980957
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_43
timestamp 1688980957
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_72
timestamp 1688980957
transform 1 0 7728 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_96
timestamp 1688980957
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_108
timestamp 1688980957
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_93
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_115
timestamp 1688980957
transform 1 0 11684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_119
timestamp 1688980957
transform 1 0 12052 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_135
timestamp 1688980957
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_145
timestamp 1688980957
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_7
timestamp 1688980957
transform 1 0 1748 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_19
timestamp 1688980957
transform 1 0 2852 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_31
timestamp 1688980957
transform 1 0 3956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_43
timestamp 1688980957
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_75
timestamp 1688980957
transform 1 0 8004 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_91
timestamp 1688980957
transform 1 0 9476 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_7
timestamp 1688980957
transform 1 0 1748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_19
timestamp 1688980957
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_105
timestamp 1688980957
transform 1 0 10764 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1688980957
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_78
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_86
timestamp 1688980957
transform 1 0 9016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_102
timestamp 1688980957
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1688980957
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_7
timestamp 1688980957
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_19
timestamp 1688980957
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_47
timestamp 1688980957
transform 1 0 5428 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_100
timestamp 1688980957
transform 1 0 10304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_104
timestamp 1688980957
transform 1 0 10672 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_126
timestamp 1688980957
transform 1 0 12696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_136
timestamp 1688980957
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_145
timestamp 1688980957
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_7
timestamp 1688980957
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_19
timestamp 1688980957
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_31
timestamp 1688980957
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_43
timestamp 1688980957
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_73
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_79
timestamp 1688980957
transform 1 0 8372 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_95
timestamp 1688980957
transform 1 0 9844 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_143
timestamp 1688980957
transform 1 0 14260 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_106
timestamp 1688980957
transform 1 0 10856 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_145
timestamp 1688980957
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_13
timestamp 1688980957
transform 1 0 2300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_25
timestamp 1688980957
transform 1 0 3404 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_37
timestamp 1688980957
transform 1 0 4508 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_49
timestamp 1688980957
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_89
timestamp 1688980957
transform 1 0 9292 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_107
timestamp 1688980957
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_7
timestamp 1688980957
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_22
timestamp 1688980957
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_76
timestamp 1688980957
transform 1 0 8096 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_101
timestamp 1688980957
transform 1 0 10396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_117
timestamp 1688980957
transform 1 0 11868 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_145
timestamp 1688980957
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_21
timestamp 1688980957
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_33
timestamp 1688980957
transform 1 0 4140 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_82
timestamp 1688980957
transform 1 0 8648 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_94
timestamp 1688980957
transform 1 0 9752 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_134
timestamp 1688980957
transform 1 0 13432 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_142
timestamp 1688980957
transform 1 0 14168 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_7
timestamp 1688980957
transform 1 0 1748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_19
timestamp 1688980957
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_100
timestamp 1688980957
transform 1 0 10304 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_104
timestamp 1688980957
transform 1 0 10672 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_123
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_145
timestamp 1688980957
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_7
timestamp 1688980957
transform 1 0 1748 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_19
timestamp 1688980957
transform 1 0 2852 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_31
timestamp 1688980957
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_43
timestamp 1688980957
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_65
timestamp 1688980957
transform 1 0 7084 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_103
timestamp 1688980957
transform 1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_72
timestamp 1688980957
transform 1 0 7728 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_145
timestamp 1688980957
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_7
timestamp 1688980957
transform 1 0 1748 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_19
timestamp 1688980957
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_31
timestamp 1688980957
transform 1 0 3956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_43
timestamp 1688980957
transform 1 0 5060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_96
timestamp 1688980957
transform 1 0 9936 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_134
timestamp 1688980957
transform 1 0 13432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_144
timestamp 1688980957
transform 1 0 14352 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_7
timestamp 1688980957
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_19
timestamp 1688980957
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_130
timestamp 1688980957
transform 1 0 13064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_145
timestamp 1688980957
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_61
timestamp 1688980957
transform 1 0 6716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_98
timestamp 1688980957
transform 1 0 10120 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_132
timestamp 1688980957
transform 1 0 13248 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_7
timestamp 1688980957
transform 1 0 1748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_19
timestamp 1688980957
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_81
timestamp 1688980957
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_105
timestamp 1688980957
transform 1 0 10764 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_145
timestamp 1688980957
transform 1 0 14444 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_7
timestamp 1688980957
transform 1 0 1748 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_19
timestamp 1688980957
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_31
timestamp 1688980957
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_43
timestamp 1688980957
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_110
timestamp 1688980957
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_88
timestamp 1688980957
transform 1 0 9200 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_100
timestamp 1688980957
transform 1 0 10304 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_111
timestamp 1688980957
transform 1 0 11316 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_144
timestamp 1688980957
transform 1 0 14352 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_7
timestamp 1688980957
transform 1 0 1748 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_13
timestamp 1688980957
transform 1 0 2300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_25
timestamp 1688980957
transform 1 0 3404 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_37
timestamp 1688980957
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_49
timestamp 1688980957
transform 1 0 5612 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_63
timestamp 1688980957
transform 1 0 6900 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_94
timestamp 1688980957
transform 1 0 9752 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_7
timestamp 1688980957
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_19
timestamp 1688980957
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_94
timestamp 1688980957
transform 1 0 9752 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_99
timestamp 1688980957
transform 1 0 10212 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_105
timestamp 1688980957
transform 1 0 10764 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_144
timestamp 1688980957
transform 1 0 14352 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_132
timestamp 1688980957
transform 1 0 13248 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_7
timestamp 1688980957
transform 1 0 1748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_19
timestamp 1688980957
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_138
timestamp 1688980957
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_144
timestamp 1688980957
transform 1 0 14352 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_7
timestamp 1688980957
transform 1 0 1748 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_19
timestamp 1688980957
transform 1 0 2852 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_31
timestamp 1688980957
transform 1 0 3956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_43
timestamp 1688980957
transform 1 0 5060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_110
timestamp 1688980957
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_8
timestamp 1688980957
transform 1 0 1840 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_20
timestamp 1688980957
transform 1 0 2944 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_92
timestamp 1688980957
transform 1 0 9568 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_104
timestamp 1688980957
transform 1 0 10672 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_144
timestamp 1688980957
transform 1 0 14352 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_10
timestamp 1688980957
transform 1 0 2024 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_22
timestamp 1688980957
transform 1 0 3128 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_34
timestamp 1688980957
transform 1 0 4232 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_46
timestamp 1688980957
transform 1 0 5336 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_54
timestamp 1688980957
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_77
timestamp 1688980957
transform 1 0 8188 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_82
timestamp 1688980957
transform 1 0 8648 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_94
timestamp 1688980957
transform 1 0 9752 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_101
timestamp 1688980957
transform 1 0 10396 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_9
timestamp 1688980957
transform 1 0 1932 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_21
timestamp 1688980957
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_90
timestamp 1688980957
transform 1 0 9384 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_102
timestamp 1688980957
transform 1 0 10488 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_110
timestamp 1688980957
transform 1 0 11224 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_129
timestamp 1688980957
transform 1 0 12972 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_136
timestamp 1688980957
transform 1 0 13616 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_9
timestamp 1688980957
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_21
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_108
timestamp 1688980957
transform 1 0 11040 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_120
timestamp 1688980957
transform 1 0 12144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_7
timestamp 1688980957
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_19
timestamp 1688980957
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_31
timestamp 1688980957
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_43
timestamp 1688980957
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_119
timestamp 1688980957
transform 1 0 12052 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_135
timestamp 1688980957
transform 1 0 13524 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_7
timestamp 1688980957
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_19
timestamp 1688980957
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_31
timestamp 1688980957
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_43
timestamp 1688980957
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_144
timestamp 1688980957
transform 1 0 14352 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_7
timestamp 1688980957
transform 1 0 1748 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_19
timestamp 1688980957
transform 1 0 2852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_88
timestamp 1688980957
transform 1 0 9200 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_94
timestamp 1688980957
transform 1 0 9752 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_106
timestamp 1688980957
transform 1 0 10856 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_118
timestamp 1688980957
transform 1 0 11960 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_132
timestamp 1688980957
transform 1 0 13248 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_87
timestamp 1688980957
transform 1 0 9108 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_91
timestamp 1688980957
transform 1 0 9476 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_100
timestamp 1688980957
transform 1 0 10304 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_131
timestamp 1688980957
transform 1 0 13156 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_144
timestamp 1688980957
transform 1 0 14352 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_7
timestamp 1688980957
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_19
timestamp 1688980957
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_145
timestamp 1688980957
transform 1 0 14444 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_7
timestamp 1688980957
transform 1 0 1748 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_19
timestamp 1688980957
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_31
timestamp 1688980957
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_43
timestamp 1688980957
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_145
timestamp 1688980957
transform 1 0 14444 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_145
timestamp 1688980957
transform 1 0 14444 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_9
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_13
timestamp 1688980957
transform 1 0 2300 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_25
timestamp 1688980957
transform 1 0 3404 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_31
timestamp 1688980957
transform 1 0 3956 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_35
timestamp 1688980957
transform 1 0 4324 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_44
timestamp 1688980957
transform 1 0 5152 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_23
timestamp 1688980957
transform 1 0 3220 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_36
timestamp 1688980957
transform 1 0 4416 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_40
timestamp 1688980957
transform 1 0 4784 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_44
timestamp 1688980957
transform 1 0 5152 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_48
timestamp 1688980957
transform 1 0 5520 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_52
timestamp 1688980957
transform 1 0 5888 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_56
timestamp 1688980957
transform 1 0 6256 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_60
timestamp 1688980957
transform 1 0 6624 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_64
timestamp 1688980957
transform 1 0 6992 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_68
timestamp 1688980957
transform 1 0 7360 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_72
timestamp 1688980957
transform 1 0 7728 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_76
timestamp 1688980957
transform 1 0 8096 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_80
timestamp 1688980957
transform 1 0 8464 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_91
timestamp 1688980957
transform 1 0 9476 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_95
timestamp 1688980957
transform 1 0 9844 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_100
timestamp 1688980957
transform 1 0 10304 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_104
timestamp 1688980957
transform 1 0 10672 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_108
timestamp 1688980957
transform 1 0 11040 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_112
timestamp 1688980957
transform 1 0 11408 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_116
timestamp 1688980957
transform 1 0 11776 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_120
timestamp 1688980957
transform 1 0 12144 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_124
timestamp 1688980957
transform 1 0 12512 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_128
timestamp 1688980957
transform 1 0 12880 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_132
timestamp 1688980957
transform 1 0 13248 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_144
timestamp 1688980957
transform 1 0 14352 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_9
timestamp 1688980957
transform 1 0 1932 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_26
timestamp 1688980957
transform 1 0 3496 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_33
timestamp 1688980957
transform 1 0 4140 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_41
timestamp 1688980957
transform 1 0 4876 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_47
timestamp 1688980957
transform 1 0 5428 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_65
timestamp 1688980957
transform 1 0 7084 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_71
timestamp 1688980957
transform 1 0 7636 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_81
timestamp 1688980957
transform 1 0 8556 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_89
timestamp 1688980957
transform 1 0 9292 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_97
timestamp 1688980957
transform 1 0 10028 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_103
timestamp 1688980957
transform 1 0 10580 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_129
timestamp 1688980957
transform 1 0 12972 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_144
timestamp 1688980957
transform 1 0 14352 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  input35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 9476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 10212 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 10948 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 11684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 12420 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input46
timestamp 1688980957
transform 1 0 2116 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input47
timestamp 1688980957
transform 1 0 2852 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  input48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1688980957
transform 1 0 4324 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1688980957
transform 1 0 5060 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 5796 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 6532 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 7268 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1688980957
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1688980957
transform 1 0 14168 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1688980957
transform 1 0 10672 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform 1 0 12420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 11776 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1688980957
transform 1 0 13616 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1688980957
transform 1 0 14168 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1688980957
transform 1 0 14168 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1688980957
transform 1 0 13616 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1688980957
transform 1 0 14168 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1688980957
transform 1 0 13064 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1688980957
transform 1 0 13616 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1688980957
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1688980957
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1688980957
transform 1 0 13248 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1688980957
transform 1 0 14168 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1688980957
transform 1 0 11684 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1688980957
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1688980957
transform 1 0 11408 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1688980957
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1688980957
transform 1 0 13064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1688980957
transform 1 0 14168 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1688980957
transform 1 0 14168 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1688980957
transform 1 0 14168 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1688980957
transform 1 0 14168 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1688980957
transform 1 0 13616 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1688980957
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1688980957
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1688980957
transform 1 0 14260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1688980957
transform 1 0 14260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input94
timestamp 1688980957
transform 1 0 11684 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1688980957
transform 1 0 13432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1688980957
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 1688980957
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1688980957
transform 1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input101
timestamp 1688980957
transform 1 0 12788 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access__0_
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access__1_
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access__2_
timestamp 1688980957
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access__3_
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_A_IO_1_bidirectional_frame_config_pass__0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_A_IO_1_bidirectional_frame_config_pass__1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_IO_1_bidirectional_frame_config_pass__2_
timestamp 1688980957
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_A_IO_1_bidirectional_frame_config_pass__3_
timestamp 1688980957
transform 1 0 5060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access__0_
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access__1_
timestamp 1688980957
transform 1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access__2_
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access__3_
timestamp 1688980957
transform 1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_B_IO_1_bidirectional_frame_config_pass__0_
timestamp 1688980957
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_B_IO_1_bidirectional_frame_config_pass__1_
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_IO_1_bidirectional_frame_config_pass__2_
timestamp 1688980957
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_B_IO_1_bidirectional_frame_config_pass__3_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit1
timestamp 1688980957
transform 1 0 10948 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit2
timestamp 1688980957
transform 1 0 6440 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit3
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit4
timestamp 1688980957
transform 1 0 10304 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit5
timestamp 1688980957
transform 1 0 11684 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit6
timestamp 1688980957
transform 1 0 6808 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit7
timestamp 1688980957
transform 1 0 8372 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit8
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit9
timestamp 1688980957
transform 1 0 11868 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit10
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit11
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit12
timestamp 1688980957
transform 1 0 10028 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit13
timestamp 1688980957
transform 1 0 12144 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit14
timestamp 1688980957
transform 1 0 7176 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit15
timestamp 1688980957
transform 1 0 6992 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit16
timestamp 1688980957
transform 1 0 10764 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit17
timestamp 1688980957
transform 1 0 11500 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit18
timestamp 1688980957
transform 1 0 8096 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit19
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit20
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit21
timestamp 1688980957
transform 1 0 11592 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit22
timestamp 1688980957
transform 1 0 6808 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit23
timestamp 1688980957
transform 1 0 7452 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit24
timestamp 1688980957
transform 1 0 5152 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit25
timestamp 1688980957
transform 1 0 8096 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit26
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit27
timestamp 1688980957
transform 1 0 10580 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit28
timestamp 1688980957
transform 1 0 10856 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit29
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit30
timestamp 1688980957
transform 1 0 6532 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit31
timestamp 1688980957
transform 1 0 5244 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit0
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit1
timestamp 1688980957
transform 1 0 9292 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit2
timestamp 1688980957
transform 1 0 7544 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit3
timestamp 1688980957
transform 1 0 9016 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit4
timestamp 1688980957
transform 1 0 12880 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit5
timestamp 1688980957
transform 1 0 12604 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit6
timestamp 1688980957
transform 1 0 7912 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit7
timestamp 1688980957
transform 1 0 9568 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit8
timestamp 1688980957
transform 1 0 12880 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit9
timestamp 1688980957
transform 1 0 12972 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit10
timestamp 1688980957
transform 1 0 11960 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit11
timestamp 1688980957
transform 1 0 12604 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit12
timestamp 1688980957
transform 1 0 4876 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit13
timestamp 1688980957
transform 1 0 6716 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit14
timestamp 1688980957
transform 1 0 9936 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit15
timestamp 1688980957
transform 1 0 10488 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit16
timestamp 1688980957
transform 1 0 11776 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit17
timestamp 1688980957
transform 1 0 13156 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit18
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit19
timestamp 1688980957
transform 1 0 6348 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit20
timestamp 1688980957
transform 1 0 7268 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit21
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit22
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit23
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit24
timestamp 1688980957
transform 1 0 12328 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit25
timestamp 1688980957
transform 1 0 12880 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit26
timestamp 1688980957
transform 1 0 7452 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit27
timestamp 1688980957
transform 1 0 8464 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit28
timestamp 1688980957
transform 1 0 11868 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit29
timestamp 1688980957
transform 1 0 10028 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit30
timestamp 1688980957
transform 1 0 7360 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit31
timestamp 1688980957
transform 1 0 8096 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit0
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit1
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit2
timestamp 1688980957
transform 1 0 9752 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit3
timestamp 1688980957
transform 1 0 10304 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit4
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit5
timestamp 1688980957
transform 1 0 11408 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit6
timestamp 1688980957
transform 1 0 7452 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit7
timestamp 1688980957
transform 1 0 8188 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit8
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit9
timestamp 1688980957
transform 1 0 11592 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit10
timestamp 1688980957
transform 1 0 12144 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit11
timestamp 1688980957
transform 1 0 12604 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit12
timestamp 1688980957
transform 1 0 9108 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit13
timestamp 1688980957
transform 1 0 9568 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit14
timestamp 1688980957
transform 1 0 5428 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit15
timestamp 1688980957
transform 1 0 5796 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit16
timestamp 1688980957
transform 1 0 12144 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit17
timestamp 1688980957
transform 1 0 12696 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit18
timestamp 1688980957
transform 1 0 6072 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit19
timestamp 1688980957
transform 1 0 7176 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit20
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit21
timestamp 1688980957
transform 1 0 12788 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit22
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit23
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit24
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit25
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit26
timestamp 1688980957
transform 1 0 10028 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit27
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit28
timestamp 1688980957
transform 1 0 12328 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit29
timestamp 1688980957
transform 1 0 12880 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit30
timestamp 1688980957
transform 1 0 4876 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit31
timestamp 1688980957
transform 1 0 5520 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit14
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit15
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit16
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit17
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit18
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit19
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit20
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit21
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit22
timestamp 1688980957
transform 1 0 9844 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit23
timestamp 1688980957
transform 1 0 5428 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit24
timestamp 1688980957
transform 1 0 5796 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit25
timestamp 1688980957
transform 1 0 9752 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit26
timestamp 1688980957
transform 1 0 6164 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit27
timestamp 1688980957
transform 1 0 6716 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit28
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit29
timestamp 1688980957
transform 1 0 9384 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit30
timestamp 1688980957
transform 1 0 7176 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit31
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__2_
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 11224 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__2_
timestamp 1688980957
transform 1 0 7544 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__3_
timestamp 1688980957
transform 1 0 6808 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__4_
timestamp 1688980957
transform 1 0 6808 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 7268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__2_
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__3_
timestamp 1688980957
transform 1 0 7268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__4_
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 7176 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 6992 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__2_
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__3_
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__4_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 11040 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 11224 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG1
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG2
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG3
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG4
timestamp 1688980957
transform 1 0 10396 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG5
timestamp 1688980957
transform 1 0 11500 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG6
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG7
timestamp 1688980957
transform 1 0 11868 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb0
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb1
timestamp 1688980957
transform 1 0 9752 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb3
timestamp 1688980957
transform 1 0 12052 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb4
timestamp 1688980957
transform 1 0 6900 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb5
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb6
timestamp 1688980957
transform 1 0 8832 0 -1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb7
timestamp 1688980957
transform 1 0 12052 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG0
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG1
timestamp 1688980957
transform 1 0 12052 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG2
timestamp 1688980957
transform 1 0 8004 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG3
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG4
timestamp 1688980957
transform 1 0 6900 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG5
timestamp 1688980957
transform -1 0 13432 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG6
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG7
timestamp 1688980957
transform 1 0 11960 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG8
timestamp 1688980957
transform 1 0 6348 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG9
timestamp 1688980957
transform 1 0 12052 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG10
timestamp 1688980957
transform 1 0 8004 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG11
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG0
timestamp 1688980957
transform 1 0 10764 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG1
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG2
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG3
timestamp 1688980957
transform 1 0 9200 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG4
timestamp 1688980957
transform 1 0 8924 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG5
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG6
timestamp 1688980957
transform 1 0 9936 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG7
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG8
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG9
timestamp 1688980957
transform 1 0 6716 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG10
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG11
timestamp 1688980957
transform 1 0 12052 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG12
timestamp 1688980957
transform 1 0 6256 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG13
timestamp 1688980957
transform 1 0 8648 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG14
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG15
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 6440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 6532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6900 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1_216 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1_218
timestamp 1688980957
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 6900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 7820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 7544 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1_217
timestamp 1688980957
transform 1 0 8464 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1_219
timestamp 1688980957
transform 1 0 6624 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6532 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 9200 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst2
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst3
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst4
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9476 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst2
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst3
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst4
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 13432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 11960 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 12052 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 11500 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 11592 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1688980957
transform 1 0 14168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 12052 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 11500 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 10948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 11500 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 13616 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 13432 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1688980957
transform 1 0 14168 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 13984 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 12052 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 13432 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 11776 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 13984 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 13432 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 10304 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 13432 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 10948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 11408 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 12880 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 13984 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output147
timestamp 1688980957
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output148
timestamp 1688980957
transform 1 0 11500 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output149
timestamp 1688980957
transform 1 0 11316 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output150
timestamp 1688980957
transform 1 0 11868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output151
timestamp 1688980957
transform 1 0 11500 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output152
timestamp 1688980957
transform 1 0 13432 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output153
timestamp 1688980957
transform 1 0 13984 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output154
timestamp 1688980957
transform 1 0 13064 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output155
timestamp 1688980957
transform 1 0 11408 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output156
timestamp 1688980957
transform 1 0 13616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output157
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output158
timestamp 1688980957
transform 1 0 10764 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output159
timestamp 1688980957
transform 1 0 13984 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output160
timestamp 1688980957
transform 1 0 12052 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output161
timestamp 1688980957
transform 1 0 13984 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output162
timestamp 1688980957
transform 1 0 13800 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output163
timestamp 1688980957
transform 1 0 12880 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output164
timestamp 1688980957
transform 1 0 12880 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output165
timestamp 1688980957
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output166
timestamp 1688980957
transform 1 0 13432 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output167
timestamp 1688980957
transform 1 0 12328 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output168
timestamp 1688980957
transform 1 0 12880 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output169
timestamp 1688980957
transform 1 0 12880 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output170
timestamp 1688980957
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1688980957
transform 1 0 14168 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output172
timestamp 1688980957
transform 1 0 13064 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1688980957
transform 1 0 14168 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output174
timestamp 1688980957
transform 1 0 13984 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output175
timestamp 1688980957
transform 1 0 13432 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output176
timestamp 1688980957
transform 1 0 13984 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output177
timestamp 1688980957
transform 1 0 12880 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1688980957
transform 1 0 14168 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1688980957
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output180
timestamp 1688980957
transform 1 0 13248 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output181
timestamp 1688980957
transform 1 0 13800 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1688980957
transform 1 0 14168 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output183
timestamp 1688980957
transform 1 0 13432 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output184
timestamp 1688980957
transform 1 0 13248 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output185
timestamp 1688980957
transform 1 0 13432 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output186
timestamp 1688980957
transform 1 0 13800 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output187
timestamp 1688980957
transform 1 0 13432 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output188
timestamp 1688980957
transform 1 0 12328 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output189
timestamp 1688980957
transform 1 0 12328 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output190
timestamp 1688980957
transform 1 0 12880 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output191
timestamp 1688980957
transform 1 0 13984 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 13432 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output193
timestamp 1688980957
transform 1 0 13432 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output194
timestamp 1688980957
transform 1 0 11776 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output195
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output197
timestamp 1688980957
transform 1 0 9476 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1688980957
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output199
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1688980957
transform 1 0 12052 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output201
timestamp 1688980957
transform 1 0 12420 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1688980957
transform 1 0 13064 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output203
timestamp 1688980957
transform 1 0 13984 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output204
timestamp 1688980957
transform 1 0 13432 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 13432 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1688980957
transform 1 0 2116 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output207
timestamp 1688980957
transform 1 0 2668 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output209
timestamp 1688980957
transform 1 0 4324 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1688980957
transform 1 0 5060 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output211
timestamp 1688980957
transform 1 0 5704 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output212
timestamp 1688980957
transform 1 0 6532 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1688980957
transform 1 0 7268 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output214
timestamp 1688980957
transform 1 0 8004 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output215
timestamp 1688980957
transform 1 0 3220 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 14812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 14812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 14812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 14812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 14812 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 14812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 14812 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 14812 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 14812 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 14812 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 14812 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 14812 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 14812 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 14812 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 14812 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 14812 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 14812 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 14812 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 14812 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 14812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 14812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 14812 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 14812 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 14812 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 14812 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 14812 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 14812 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 14812 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 14812 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 14812 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 14812 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 14812 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 14812 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 14812 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 1564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 2024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 3128 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 4048 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 4876 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 5612 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 7084 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 7820 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 8464 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 10028 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 12236 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 12880 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 13984 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 1748 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 2024 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 2760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 3312 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 4140 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 5612 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 6348 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 7084 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 7820 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 8556 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 9200 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform -1 0 10304 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 10764 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 11500 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 12236 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 12972 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 11432 160 11552 0 FreeSans 480 0 0 0 A_I_top
port 0 nsew signal tristate
flabel metal3 s 0 9800 160 9920 0 FreeSans 480 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s 0 10616 160 10736 0 FreeSans 480 0 0 0 A_T_top
port 2 nsew signal tristate
flabel metal3 s 0 12248 160 12368 0 FreeSans 480 0 0 0 A_config_C_bit0
port 3 nsew signal tristate
flabel metal3 s 0 13064 160 13184 0 FreeSans 480 0 0 0 A_config_C_bit1
port 4 nsew signal tristate
flabel metal3 s 0 13880 160 14000 0 FreeSans 480 0 0 0 A_config_C_bit2
port 5 nsew signal tristate
flabel metal3 s 0 14696 160 14816 0 FreeSans 480 0 0 0 A_config_C_bit3
port 6 nsew signal tristate
flabel metal3 s 0 5720 160 5840 0 FreeSans 480 0 0 0 B_I_top
port 7 nsew signal tristate
flabel metal3 s 0 4088 160 4208 0 FreeSans 480 0 0 0 B_O_top
port 8 nsew signal input
flabel metal3 s 0 4904 160 5024 0 FreeSans 480 0 0 0 B_T_top
port 9 nsew signal tristate
flabel metal3 s 0 6536 160 6656 0 FreeSans 480 0 0 0 B_config_C_bit0
port 10 nsew signal tristate
flabel metal3 s 0 7352 160 7472 0 FreeSans 480 0 0 0 B_config_C_bit1
port 11 nsew signal tristate
flabel metal3 s 0 8168 160 8288 0 FreeSans 480 0 0 0 B_config_C_bit2
port 12 nsew signal tristate
flabel metal3 s 0 8984 160 9104 0 FreeSans 480 0 0 0 B_config_C_bit3
port 13 nsew signal tristate
flabel metal3 s 15840 18232 16000 18352 0 FreeSans 480 0 0 0 E1BEG[0]
port 14 nsew signal tristate
flabel metal3 s 15840 18504 16000 18624 0 FreeSans 480 0 0 0 E1BEG[1]
port 15 nsew signal tristate
flabel metal3 s 15840 18776 16000 18896 0 FreeSans 480 0 0 0 E1BEG[2]
port 16 nsew signal tristate
flabel metal3 s 15840 19048 16000 19168 0 FreeSans 480 0 0 0 E1BEG[3]
port 17 nsew signal tristate
flabel metal3 s 15840 19320 16000 19440 0 FreeSans 480 0 0 0 E2BEG[0]
port 18 nsew signal tristate
flabel metal3 s 15840 19592 16000 19712 0 FreeSans 480 0 0 0 E2BEG[1]
port 19 nsew signal tristate
flabel metal3 s 15840 19864 16000 19984 0 FreeSans 480 0 0 0 E2BEG[2]
port 20 nsew signal tristate
flabel metal3 s 15840 20136 16000 20256 0 FreeSans 480 0 0 0 E2BEG[3]
port 21 nsew signal tristate
flabel metal3 s 15840 20408 16000 20528 0 FreeSans 480 0 0 0 E2BEG[4]
port 22 nsew signal tristate
flabel metal3 s 15840 20680 16000 20800 0 FreeSans 480 0 0 0 E2BEG[5]
port 23 nsew signal tristate
flabel metal3 s 15840 20952 16000 21072 0 FreeSans 480 0 0 0 E2BEG[6]
port 24 nsew signal tristate
flabel metal3 s 15840 21224 16000 21344 0 FreeSans 480 0 0 0 E2BEG[7]
port 25 nsew signal tristate
flabel metal3 s 15840 21496 16000 21616 0 FreeSans 480 0 0 0 E2BEGb[0]
port 26 nsew signal tristate
flabel metal3 s 15840 21768 16000 21888 0 FreeSans 480 0 0 0 E2BEGb[1]
port 27 nsew signal tristate
flabel metal3 s 15840 22040 16000 22160 0 FreeSans 480 0 0 0 E2BEGb[2]
port 28 nsew signal tristate
flabel metal3 s 15840 22312 16000 22432 0 FreeSans 480 0 0 0 E2BEGb[3]
port 29 nsew signal tristate
flabel metal3 s 15840 22584 16000 22704 0 FreeSans 480 0 0 0 E2BEGb[4]
port 30 nsew signal tristate
flabel metal3 s 15840 22856 16000 22976 0 FreeSans 480 0 0 0 E2BEGb[5]
port 31 nsew signal tristate
flabel metal3 s 15840 23128 16000 23248 0 FreeSans 480 0 0 0 E2BEGb[6]
port 32 nsew signal tristate
flabel metal3 s 15840 23400 16000 23520 0 FreeSans 480 0 0 0 E2BEGb[7]
port 33 nsew signal tristate
flabel metal3 s 15840 28024 16000 28144 0 FreeSans 480 0 0 0 E6BEG[0]
port 34 nsew signal tristate
flabel metal3 s 15840 30744 16000 30864 0 FreeSans 480 0 0 0 E6BEG[10]
port 35 nsew signal tristate
flabel metal3 s 15840 31016 16000 31136 0 FreeSans 480 0 0 0 E6BEG[11]
port 36 nsew signal tristate
flabel metal3 s 15840 28296 16000 28416 0 FreeSans 480 0 0 0 E6BEG[1]
port 37 nsew signal tristate
flabel metal3 s 15840 28568 16000 28688 0 FreeSans 480 0 0 0 E6BEG[2]
port 38 nsew signal tristate
flabel metal3 s 15840 28840 16000 28960 0 FreeSans 480 0 0 0 E6BEG[3]
port 39 nsew signal tristate
flabel metal3 s 15840 29112 16000 29232 0 FreeSans 480 0 0 0 E6BEG[4]
port 40 nsew signal tristate
flabel metal3 s 15840 29384 16000 29504 0 FreeSans 480 0 0 0 E6BEG[5]
port 41 nsew signal tristate
flabel metal3 s 15840 29656 16000 29776 0 FreeSans 480 0 0 0 E6BEG[6]
port 42 nsew signal tristate
flabel metal3 s 15840 29928 16000 30048 0 FreeSans 480 0 0 0 E6BEG[7]
port 43 nsew signal tristate
flabel metal3 s 15840 30200 16000 30320 0 FreeSans 480 0 0 0 E6BEG[8]
port 44 nsew signal tristate
flabel metal3 s 15840 30472 16000 30592 0 FreeSans 480 0 0 0 E6BEG[9]
port 45 nsew signal tristate
flabel metal3 s 15840 23672 16000 23792 0 FreeSans 480 0 0 0 EE4BEG[0]
port 46 nsew signal tristate
flabel metal3 s 15840 26392 16000 26512 0 FreeSans 480 0 0 0 EE4BEG[10]
port 47 nsew signal tristate
flabel metal3 s 15840 26664 16000 26784 0 FreeSans 480 0 0 0 EE4BEG[11]
port 48 nsew signal tristate
flabel metal3 s 15840 26936 16000 27056 0 FreeSans 480 0 0 0 EE4BEG[12]
port 49 nsew signal tristate
flabel metal3 s 15840 27208 16000 27328 0 FreeSans 480 0 0 0 EE4BEG[13]
port 50 nsew signal tristate
flabel metal3 s 15840 27480 16000 27600 0 FreeSans 480 0 0 0 EE4BEG[14]
port 51 nsew signal tristate
flabel metal3 s 15840 27752 16000 27872 0 FreeSans 480 0 0 0 EE4BEG[15]
port 52 nsew signal tristate
flabel metal3 s 15840 23944 16000 24064 0 FreeSans 480 0 0 0 EE4BEG[1]
port 53 nsew signal tristate
flabel metal3 s 15840 24216 16000 24336 0 FreeSans 480 0 0 0 EE4BEG[2]
port 54 nsew signal tristate
flabel metal3 s 15840 24488 16000 24608 0 FreeSans 480 0 0 0 EE4BEG[3]
port 55 nsew signal tristate
flabel metal3 s 15840 24760 16000 24880 0 FreeSans 480 0 0 0 EE4BEG[4]
port 56 nsew signal tristate
flabel metal3 s 15840 25032 16000 25152 0 FreeSans 480 0 0 0 EE4BEG[5]
port 57 nsew signal tristate
flabel metal3 s 15840 25304 16000 25424 0 FreeSans 480 0 0 0 EE4BEG[6]
port 58 nsew signal tristate
flabel metal3 s 15840 25576 16000 25696 0 FreeSans 480 0 0 0 EE4BEG[7]
port 59 nsew signal tristate
flabel metal3 s 15840 25848 16000 25968 0 FreeSans 480 0 0 0 EE4BEG[8]
port 60 nsew signal tristate
flabel metal3 s 15840 26120 16000 26240 0 FreeSans 480 0 0 0 EE4BEG[9]
port 61 nsew signal tristate
flabel metal3 s 0 15512 160 15632 0 FreeSans 480 0 0 0 FrameData[0]
port 62 nsew signal input
flabel metal3 s 0 23672 160 23792 0 FreeSans 480 0 0 0 FrameData[10]
port 63 nsew signal input
flabel metal3 s 0 24488 160 24608 0 FreeSans 480 0 0 0 FrameData[11]
port 64 nsew signal input
flabel metal3 s 0 25304 160 25424 0 FreeSans 480 0 0 0 FrameData[12]
port 65 nsew signal input
flabel metal3 s 0 26120 160 26240 0 FreeSans 480 0 0 0 FrameData[13]
port 66 nsew signal input
flabel metal3 s 0 26936 160 27056 0 FreeSans 480 0 0 0 FrameData[14]
port 67 nsew signal input
flabel metal3 s 0 27752 160 27872 0 FreeSans 480 0 0 0 FrameData[15]
port 68 nsew signal input
flabel metal3 s 0 28568 160 28688 0 FreeSans 480 0 0 0 FrameData[16]
port 69 nsew signal input
flabel metal3 s 0 29384 160 29504 0 FreeSans 480 0 0 0 FrameData[17]
port 70 nsew signal input
flabel metal3 s 0 30200 160 30320 0 FreeSans 480 0 0 0 FrameData[18]
port 71 nsew signal input
flabel metal3 s 0 31016 160 31136 0 FreeSans 480 0 0 0 FrameData[19]
port 72 nsew signal input
flabel metal3 s 0 16328 160 16448 0 FreeSans 480 0 0 0 FrameData[1]
port 73 nsew signal input
flabel metal3 s 0 31832 160 31952 0 FreeSans 480 0 0 0 FrameData[20]
port 74 nsew signal input
flabel metal3 s 0 32648 160 32768 0 FreeSans 480 0 0 0 FrameData[21]
port 75 nsew signal input
flabel metal3 s 0 33464 160 33584 0 FreeSans 480 0 0 0 FrameData[22]
port 76 nsew signal input
flabel metal3 s 0 34280 160 34400 0 FreeSans 480 0 0 0 FrameData[23]
port 77 nsew signal input
flabel metal3 s 0 35096 160 35216 0 FreeSans 480 0 0 0 FrameData[24]
port 78 nsew signal input
flabel metal3 s 0 35912 160 36032 0 FreeSans 480 0 0 0 FrameData[25]
port 79 nsew signal input
flabel metal3 s 0 36728 160 36848 0 FreeSans 480 0 0 0 FrameData[26]
port 80 nsew signal input
flabel metal3 s 0 37544 160 37664 0 FreeSans 480 0 0 0 FrameData[27]
port 81 nsew signal input
flabel metal3 s 0 38360 160 38480 0 FreeSans 480 0 0 0 FrameData[28]
port 82 nsew signal input
flabel metal3 s 0 39176 160 39296 0 FreeSans 480 0 0 0 FrameData[29]
port 83 nsew signal input
flabel metal3 s 0 17144 160 17264 0 FreeSans 480 0 0 0 FrameData[2]
port 84 nsew signal input
flabel metal3 s 0 39992 160 40112 0 FreeSans 480 0 0 0 FrameData[30]
port 85 nsew signal input
flabel metal3 s 0 40808 160 40928 0 FreeSans 480 0 0 0 FrameData[31]
port 86 nsew signal input
flabel metal3 s 0 17960 160 18080 0 FreeSans 480 0 0 0 FrameData[3]
port 87 nsew signal input
flabel metal3 s 0 18776 160 18896 0 FreeSans 480 0 0 0 FrameData[4]
port 88 nsew signal input
flabel metal3 s 0 19592 160 19712 0 FreeSans 480 0 0 0 FrameData[5]
port 89 nsew signal input
flabel metal3 s 0 20408 160 20528 0 FreeSans 480 0 0 0 FrameData[6]
port 90 nsew signal input
flabel metal3 s 0 21224 160 21344 0 FreeSans 480 0 0 0 FrameData[7]
port 91 nsew signal input
flabel metal3 s 0 22040 160 22160 0 FreeSans 480 0 0 0 FrameData[8]
port 92 nsew signal input
flabel metal3 s 0 22856 160 22976 0 FreeSans 480 0 0 0 FrameData[9]
port 93 nsew signal input
flabel metal3 s 15840 31288 16000 31408 0 FreeSans 480 0 0 0 FrameData_O[0]
port 94 nsew signal tristate
flabel metal3 s 15840 34008 16000 34128 0 FreeSans 480 0 0 0 FrameData_O[10]
port 95 nsew signal tristate
flabel metal3 s 15840 34280 16000 34400 0 FreeSans 480 0 0 0 FrameData_O[11]
port 96 nsew signal tristate
flabel metal3 s 15840 34552 16000 34672 0 FreeSans 480 0 0 0 FrameData_O[12]
port 97 nsew signal tristate
flabel metal3 s 15840 34824 16000 34944 0 FreeSans 480 0 0 0 FrameData_O[13]
port 98 nsew signal tristate
flabel metal3 s 15840 35096 16000 35216 0 FreeSans 480 0 0 0 FrameData_O[14]
port 99 nsew signal tristate
flabel metal3 s 15840 35368 16000 35488 0 FreeSans 480 0 0 0 FrameData_O[15]
port 100 nsew signal tristate
flabel metal3 s 15840 35640 16000 35760 0 FreeSans 480 0 0 0 FrameData_O[16]
port 101 nsew signal tristate
flabel metal3 s 15840 35912 16000 36032 0 FreeSans 480 0 0 0 FrameData_O[17]
port 102 nsew signal tristate
flabel metal3 s 15840 36184 16000 36304 0 FreeSans 480 0 0 0 FrameData_O[18]
port 103 nsew signal tristate
flabel metal3 s 15840 36456 16000 36576 0 FreeSans 480 0 0 0 FrameData_O[19]
port 104 nsew signal tristate
flabel metal3 s 15840 31560 16000 31680 0 FreeSans 480 0 0 0 FrameData_O[1]
port 105 nsew signal tristate
flabel metal3 s 15840 36728 16000 36848 0 FreeSans 480 0 0 0 FrameData_O[20]
port 106 nsew signal tristate
flabel metal3 s 15840 37000 16000 37120 0 FreeSans 480 0 0 0 FrameData_O[21]
port 107 nsew signal tristate
flabel metal3 s 15840 37272 16000 37392 0 FreeSans 480 0 0 0 FrameData_O[22]
port 108 nsew signal tristate
flabel metal3 s 15840 37544 16000 37664 0 FreeSans 480 0 0 0 FrameData_O[23]
port 109 nsew signal tristate
flabel metal3 s 15840 37816 16000 37936 0 FreeSans 480 0 0 0 FrameData_O[24]
port 110 nsew signal tristate
flabel metal3 s 15840 38088 16000 38208 0 FreeSans 480 0 0 0 FrameData_O[25]
port 111 nsew signal tristate
flabel metal3 s 15840 38360 16000 38480 0 FreeSans 480 0 0 0 FrameData_O[26]
port 112 nsew signal tristate
flabel metal3 s 15840 38632 16000 38752 0 FreeSans 480 0 0 0 FrameData_O[27]
port 113 nsew signal tristate
flabel metal3 s 15840 38904 16000 39024 0 FreeSans 480 0 0 0 FrameData_O[28]
port 114 nsew signal tristate
flabel metal3 s 15840 39176 16000 39296 0 FreeSans 480 0 0 0 FrameData_O[29]
port 115 nsew signal tristate
flabel metal3 s 15840 31832 16000 31952 0 FreeSans 480 0 0 0 FrameData_O[2]
port 116 nsew signal tristate
flabel metal3 s 15840 39448 16000 39568 0 FreeSans 480 0 0 0 FrameData_O[30]
port 117 nsew signal tristate
flabel metal3 s 15840 39720 16000 39840 0 FreeSans 480 0 0 0 FrameData_O[31]
port 118 nsew signal tristate
flabel metal3 s 15840 32104 16000 32224 0 FreeSans 480 0 0 0 FrameData_O[3]
port 119 nsew signal tristate
flabel metal3 s 15840 32376 16000 32496 0 FreeSans 480 0 0 0 FrameData_O[4]
port 120 nsew signal tristate
flabel metal3 s 15840 32648 16000 32768 0 FreeSans 480 0 0 0 FrameData_O[5]
port 121 nsew signal tristate
flabel metal3 s 15840 32920 16000 33040 0 FreeSans 480 0 0 0 FrameData_O[6]
port 122 nsew signal tristate
flabel metal3 s 15840 33192 16000 33312 0 FreeSans 480 0 0 0 FrameData_O[7]
port 123 nsew signal tristate
flabel metal3 s 15840 33464 16000 33584 0 FreeSans 480 0 0 0 FrameData_O[8]
port 124 nsew signal tristate
flabel metal3 s 15840 33736 16000 33856 0 FreeSans 480 0 0 0 FrameData_O[9]
port 125 nsew signal tristate
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 126 nsew signal input
flabel metal2 s 8666 0 8722 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 127 nsew signal input
flabel metal2 s 9402 0 9458 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 128 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 129 nsew signal input
flabel metal2 s 10874 0 10930 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 130 nsew signal input
flabel metal2 s 11610 0 11666 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 131 nsew signal input
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 132 nsew signal input
flabel metal2 s 13082 0 13138 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 133 nsew signal input
flabel metal2 s 13818 0 13874 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 134 nsew signal input
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 135 nsew signal input
flabel metal2 s 15290 0 15346 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 136 nsew signal input
flabel metal2 s 2042 0 2098 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 137 nsew signal input
flabel metal2 s 2778 0 2834 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 138 nsew signal input
flabel metal2 s 3514 0 3570 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 139 nsew signal input
flabel metal2 s 4250 0 4306 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 140 nsew signal input
flabel metal2 s 4986 0 5042 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 141 nsew signal input
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 142 nsew signal input
flabel metal2 s 6458 0 6514 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 143 nsew signal input
flabel metal2 s 7194 0 7250 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 144 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 145 nsew signal input
flabel metal2 s 1306 44840 1362 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 146 nsew signal tristate
flabel metal2 s 8666 44840 8722 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 147 nsew signal tristate
flabel metal2 s 9402 44840 9458 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 148 nsew signal tristate
flabel metal2 s 10138 44840 10194 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 149 nsew signal tristate
flabel metal2 s 10874 44840 10930 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 150 nsew signal tristate
flabel metal2 s 11610 44840 11666 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 151 nsew signal tristate
flabel metal2 s 12346 44840 12402 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 152 nsew signal tristate
flabel metal2 s 13082 44840 13138 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 153 nsew signal tristate
flabel metal2 s 13818 44840 13874 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 154 nsew signal tristate
flabel metal2 s 14554 44840 14610 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 155 nsew signal tristate
flabel metal2 s 15290 44840 15346 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 156 nsew signal tristate
flabel metal2 s 2042 44840 2098 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 157 nsew signal tristate
flabel metal2 s 2778 44840 2834 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 158 nsew signal tristate
flabel metal2 s 3514 44840 3570 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 159 nsew signal tristate
flabel metal2 s 4250 44840 4306 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 160 nsew signal tristate
flabel metal2 s 4986 44840 5042 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 161 nsew signal tristate
flabel metal2 s 5722 44840 5778 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 162 nsew signal tristate
flabel metal2 s 6458 44840 6514 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 163 nsew signal tristate
flabel metal2 s 7194 44840 7250 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 164 nsew signal tristate
flabel metal2 s 7930 44840 7986 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 165 nsew signal tristate
flabel metal2 s 570 0 626 160 0 FreeSans 224 90 0 0 UserCLK
port 166 nsew signal input
flabel metal2 s 570 44840 626 45000 0 FreeSans 224 90 0 0 UserCLKo
port 167 nsew signal tristate
flabel metal4 s 4370 1040 4690 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 7797 1040 8117 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 11224 1040 11544 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 14651 1040 14971 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 2657 1040 2977 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 6084 1040 6404 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 9511 1040 9831 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 12938 1040 13258 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal3 s 15840 5176 16000 5296 0 FreeSans 480 0 0 0 W1END[0]
port 170 nsew signal input
flabel metal3 s 15840 5448 16000 5568 0 FreeSans 480 0 0 0 W1END[1]
port 171 nsew signal input
flabel metal3 s 15840 5720 16000 5840 0 FreeSans 480 0 0 0 W1END[2]
port 172 nsew signal input
flabel metal3 s 15840 5992 16000 6112 0 FreeSans 480 0 0 0 W1END[3]
port 173 nsew signal input
flabel metal3 s 15840 8440 16000 8560 0 FreeSans 480 0 0 0 W2END[0]
port 174 nsew signal input
flabel metal3 s 15840 8712 16000 8832 0 FreeSans 480 0 0 0 W2END[1]
port 175 nsew signal input
flabel metal3 s 15840 8984 16000 9104 0 FreeSans 480 0 0 0 W2END[2]
port 176 nsew signal input
flabel metal3 s 15840 9256 16000 9376 0 FreeSans 480 0 0 0 W2END[3]
port 177 nsew signal input
flabel metal3 s 15840 9528 16000 9648 0 FreeSans 480 0 0 0 W2END[4]
port 178 nsew signal input
flabel metal3 s 15840 9800 16000 9920 0 FreeSans 480 0 0 0 W2END[5]
port 179 nsew signal input
flabel metal3 s 15840 10072 16000 10192 0 FreeSans 480 0 0 0 W2END[6]
port 180 nsew signal input
flabel metal3 s 15840 10344 16000 10464 0 FreeSans 480 0 0 0 W2END[7]
port 181 nsew signal input
flabel metal3 s 15840 6264 16000 6384 0 FreeSans 480 0 0 0 W2MID[0]
port 182 nsew signal input
flabel metal3 s 15840 6536 16000 6656 0 FreeSans 480 0 0 0 W2MID[1]
port 183 nsew signal input
flabel metal3 s 15840 6808 16000 6928 0 FreeSans 480 0 0 0 W2MID[2]
port 184 nsew signal input
flabel metal3 s 15840 7080 16000 7200 0 FreeSans 480 0 0 0 W2MID[3]
port 185 nsew signal input
flabel metal3 s 15840 7352 16000 7472 0 FreeSans 480 0 0 0 W2MID[4]
port 186 nsew signal input
flabel metal3 s 15840 7624 16000 7744 0 FreeSans 480 0 0 0 W2MID[5]
port 187 nsew signal input
flabel metal3 s 15840 7896 16000 8016 0 FreeSans 480 0 0 0 W2MID[6]
port 188 nsew signal input
flabel metal3 s 15840 8168 16000 8288 0 FreeSans 480 0 0 0 W2MID[7]
port 189 nsew signal input
flabel metal3 s 15840 14968 16000 15088 0 FreeSans 480 0 0 0 W6END[0]
port 190 nsew signal input
flabel metal3 s 15840 17688 16000 17808 0 FreeSans 480 0 0 0 W6END[10]
port 191 nsew signal input
flabel metal3 s 15840 17960 16000 18080 0 FreeSans 480 0 0 0 W6END[11]
port 192 nsew signal input
flabel metal3 s 15840 15240 16000 15360 0 FreeSans 480 0 0 0 W6END[1]
port 193 nsew signal input
flabel metal3 s 15840 15512 16000 15632 0 FreeSans 480 0 0 0 W6END[2]
port 194 nsew signal input
flabel metal3 s 15840 15784 16000 15904 0 FreeSans 480 0 0 0 W6END[3]
port 195 nsew signal input
flabel metal3 s 15840 16056 16000 16176 0 FreeSans 480 0 0 0 W6END[4]
port 196 nsew signal input
flabel metal3 s 15840 16328 16000 16448 0 FreeSans 480 0 0 0 W6END[5]
port 197 nsew signal input
flabel metal3 s 15840 16600 16000 16720 0 FreeSans 480 0 0 0 W6END[6]
port 198 nsew signal input
flabel metal3 s 15840 16872 16000 16992 0 FreeSans 480 0 0 0 W6END[7]
port 199 nsew signal input
flabel metal3 s 15840 17144 16000 17264 0 FreeSans 480 0 0 0 W6END[8]
port 200 nsew signal input
flabel metal3 s 15840 17416 16000 17536 0 FreeSans 480 0 0 0 W6END[9]
port 201 nsew signal input
flabel metal3 s 15840 10616 16000 10736 0 FreeSans 480 0 0 0 WW4END[0]
port 202 nsew signal input
flabel metal3 s 15840 13336 16000 13456 0 FreeSans 480 0 0 0 WW4END[10]
port 203 nsew signal input
flabel metal3 s 15840 13608 16000 13728 0 FreeSans 480 0 0 0 WW4END[11]
port 204 nsew signal input
flabel metal3 s 15840 13880 16000 14000 0 FreeSans 480 0 0 0 WW4END[12]
port 205 nsew signal input
flabel metal3 s 15840 14152 16000 14272 0 FreeSans 480 0 0 0 WW4END[13]
port 206 nsew signal input
flabel metal3 s 15840 14424 16000 14544 0 FreeSans 480 0 0 0 WW4END[14]
port 207 nsew signal input
flabel metal3 s 15840 14696 16000 14816 0 FreeSans 480 0 0 0 WW4END[15]
port 208 nsew signal input
flabel metal3 s 15840 10888 16000 11008 0 FreeSans 480 0 0 0 WW4END[1]
port 209 nsew signal input
flabel metal3 s 15840 11160 16000 11280 0 FreeSans 480 0 0 0 WW4END[2]
port 210 nsew signal input
flabel metal3 s 15840 11432 16000 11552 0 FreeSans 480 0 0 0 WW4END[3]
port 211 nsew signal input
flabel metal3 s 15840 11704 16000 11824 0 FreeSans 480 0 0 0 WW4END[4]
port 212 nsew signal input
flabel metal3 s 15840 11976 16000 12096 0 FreeSans 480 0 0 0 WW4END[5]
port 213 nsew signal input
flabel metal3 s 15840 12248 16000 12368 0 FreeSans 480 0 0 0 WW4END[6]
port 214 nsew signal input
flabel metal3 s 15840 12520 16000 12640 0 FreeSans 480 0 0 0 WW4END[7]
port 215 nsew signal input
flabel metal3 s 15840 12792 16000 12912 0 FreeSans 480 0 0 0 WW4END[8]
port 216 nsew signal input
flabel metal3 s 15840 13064 16000 13184 0 FreeSans 480 0 0 0 WW4END[9]
port 217 nsew signal input
rlabel via1 8037 43520 8037 43520 0 VGND
rlabel metal1 7958 42976 7958 42976 0 VPWR
rlabel metal1 2277 10642 2277 10642 0 A_I
rlabel metal3 498 11492 498 11492 0 A_I_top
rlabel metal1 10994 18734 10994 18734 0 A_O
rlabel metal3 590 9860 590 9860 0 A_O_top
rlabel metal1 7176 27642 7176 27642 0 A_Q
rlabel metal1 6716 9146 6716 9146 0 A_T
rlabel metal3 475 10676 475 10676 0 A_T_top
rlabel metal3 498 12308 498 12308 0 A_config_C_bit0
rlabel metal3 498 13124 498 13124 0 A_config_C_bit1
rlabel metal3 498 13940 498 13940 0 A_config_C_bit2
rlabel metal3 498 14756 498 14756 0 A_config_C_bit3
rlabel metal2 13386 5933 13386 5933 0 B_I
rlabel metal3 498 5780 498 5780 0 B_I_top
rlabel metal2 9430 21454 9430 21454 0 B_O
rlabel metal3 452 4148 452 4148 0 B_O_top
rlabel metal1 8464 20230 8464 20230 0 B_Q
rlabel metal1 2070 5712 2070 5712 0 B_T
rlabel metal3 498 4964 498 4964 0 B_T_top
rlabel metal3 498 6596 498 6596 0 B_config_C_bit0
rlabel metal3 498 7412 498 7412 0 B_config_C_bit1
rlabel metal3 912 8228 912 8228 0 B_config_C_bit2
rlabel metal3 199 9044 199 9044 0 B_config_C_bit3
rlabel metal1 2300 12206 2300 12206 0 ConfigBits\[0\]
rlabel metal1 9614 6426 9614 6426 0 ConfigBits\[100\]
rlabel metal2 10718 7446 10718 7446 0 ConfigBits\[101\]
rlabel metal1 12190 8602 12190 8602 0 ConfigBits\[102\]
rlabel metal2 12374 8500 12374 8500 0 ConfigBits\[103\]
rlabel metal1 7866 8330 7866 8330 0 ConfigBits\[104\]
rlabel metal1 8326 9010 8326 9010 0 ConfigBits\[105\]
rlabel metal1 6532 8942 6532 8942 0 ConfigBits\[106\]
rlabel metal1 10212 8330 10212 8330 0 ConfigBits\[107\]
rlabel metal2 10718 9486 10718 9486 0 ConfigBits\[108\]
rlabel metal1 11914 4794 11914 4794 0 ConfigBits\[109\]
rlabel metal1 7084 19958 7084 19958 0 ConfigBits\[10\]
rlabel metal2 12742 6086 12742 6086 0 ConfigBits\[110\]
rlabel metal1 7084 10506 7084 10506 0 ConfigBits\[111\]
rlabel metal2 7774 10710 7774 10710 0 ConfigBits\[112\]
rlabel metal1 6210 10642 6210 10642 0 ConfigBits\[113\]
rlabel metal1 10994 20434 10994 20434 0 ConfigBits\[11\]
rlabel metal1 7636 17102 7636 17102 0 ConfigBits\[12\]
rlabel metal1 8050 16762 8050 16762 0 ConfigBits\[13\]
rlabel metal1 9798 17034 9798 17034 0 ConfigBits\[14\]
rlabel metal2 10718 17340 10718 17340 0 ConfigBits\[15\]
rlabel metal1 8740 15946 8740 15946 0 ConfigBits\[16\]
rlabel metal2 9982 15844 9982 15844 0 ConfigBits\[17\]
rlabel metal2 13294 17986 13294 17986 0 ConfigBits\[18\]
rlabel metal2 13846 18428 13846 18428 0 ConfigBits\[19\]
rlabel metal1 2300 13906 2300 13906 0 ConfigBits\[1\]
rlabel metal1 11086 14552 11086 14552 0 ConfigBits\[20\]
rlabel metal2 11638 14892 11638 14892 0 ConfigBits\[21\]
rlabel metal2 12558 13600 12558 13600 0 ConfigBits\[22\]
rlabel metal1 12604 12410 12604 12410 0 ConfigBits\[23\]
rlabel metal1 9062 19958 9062 19958 0 ConfigBits\[24\]
rlabel metal2 9246 20128 9246 20128 0 ConfigBits\[25\]
rlabel metal2 12558 16422 12558 16422 0 ConfigBits\[26\]
rlabel metal2 13064 16558 13064 16558 0 ConfigBits\[27\]
rlabel metal1 13248 21862 13248 21862 0 ConfigBits\[28\]
rlabel metal1 13754 21114 13754 21114 0 ConfigBits\[29\]
rlabel metal1 2300 14994 2300 14994 0 ConfigBits\[2\]
rlabel metal1 10304 22066 10304 22066 0 ConfigBits\[30\]
rlabel metal1 10810 25670 10810 25670 0 ConfigBits\[31\]
rlabel metal2 6486 15130 6486 15130 0 ConfigBits\[32\]
rlabel metal1 6900 14586 6900 14586 0 ConfigBits\[33\]
rlabel metal1 12696 19958 12696 19958 0 ConfigBits\[34\]
rlabel metal1 13524 19482 13524 19482 0 ConfigBits\[35\]
rlabel metal1 7360 13498 7360 13498 0 ConfigBits\[36\]
rlabel metal2 8142 13974 8142 13974 0 ConfigBits\[37\]
rlabel metal1 13202 11322 13202 11322 0 ConfigBits\[38\]
rlabel metal2 13846 11254 13846 11254 0 ConfigBits\[39\]
rlabel metal1 2208 16422 2208 16422 0 ConfigBits\[3\]
rlabel metal2 8510 13668 8510 13668 0 ConfigBits\[40\]
rlabel metal1 9706 13498 9706 13498 0 ConfigBits\[41\]
rlabel metal3 13340 10132 13340 10132 0 ConfigBits\[42\]
rlabel metal1 12880 7514 12880 7514 0 ConfigBits\[43\]
rlabel metal2 11454 24446 11454 24446 0 ConfigBits\[44\]
rlabel metal2 12558 24480 12558 24480 0 ConfigBits\[45\]
rlabel metal1 13340 23290 13340 23290 0 ConfigBits\[46\]
rlabel metal2 13846 24140 13846 24140 0 ConfigBits\[47\]
rlabel metal1 6486 23562 6486 23562 0 ConfigBits\[48\]
rlabel metal2 7590 23868 7590 23868 0 ConfigBits\[49\]
rlabel metal1 2392 6426 2392 6426 0 ConfigBits\[4\]
rlabel metal1 9936 28662 9936 28662 0 ConfigBits\[50\]
rlabel metal2 10442 29852 10442 29852 0 ConfigBits\[51\]
rlabel metal1 8602 11628 8602 11628 0 ConfigBits\[52\]
rlabel metal2 10074 11560 10074 11560 0 ConfigBits\[53\]
rlabel metal2 13294 13192 13294 13192 0 ConfigBits\[54\]
rlabel metal2 13846 13532 13846 13532 0 ConfigBits\[55\]
rlabel metal1 9798 16694 9798 16694 0 ConfigBits\[56\]
rlabel metal1 10856 20230 10856 20230 0 ConfigBits\[57\]
rlabel metal1 12742 15640 12742 15640 0 ConfigBits\[58\]
rlabel metal1 13662 15130 13662 15130 0 ConfigBits\[59\]
rlabel metal1 2530 6766 2530 6766 0 ConfigBits\[5\]
rlabel metal1 13156 25466 13156 25466 0 ConfigBits\[60\]
rlabel metal2 13846 26588 13846 26588 0 ConfigBits\[61\]
rlabel metal1 6670 26826 6670 26826 0 ConfigBits\[62\]
rlabel metal1 7866 26554 7866 26554 0 ConfigBits\[63\]
rlabel metal1 11592 26826 11592 26826 0 ConfigBits\[64\]
rlabel metal2 11546 26656 11546 26656 0 ConfigBits\[65\]
rlabel metal1 12788 26486 12788 26486 0 ConfigBits\[66\]
rlabel metal1 13616 26418 13616 26418 0 ConfigBits\[67\]
rlabel metal1 6440 27574 6440 27574 0 ConfigBits\[68\]
rlabel metal1 7452 28390 7452 28390 0 ConfigBits\[69\]
rlabel metal1 2300 8466 2300 8466 0 ConfigBits\[6\]
rlabel metal1 8832 27914 8832 27914 0 ConfigBits\[70\]
rlabel metal1 9936 27642 9936 27642 0 ConfigBits\[71\]
rlabel metal2 13294 6154 13294 6154 0 ConfigBits\[72\]
rlabel metal1 13570 4794 13570 4794 0 ConfigBits\[73\]
rlabel metal1 13478 5338 13478 5338 0 ConfigBits\[74\]
rlabel metal1 13892 3910 13892 3910 0 ConfigBits\[75\]
rlabel metal1 9062 25398 9062 25398 0 ConfigBits\[76\]
rlabel metal2 9522 25126 9522 25126 0 ConfigBits\[77\]
rlabel metal1 12788 28662 12788 28662 0 ConfigBits\[78\]
rlabel metal2 11086 28849 11086 28849 0 ConfigBits\[79\]
rlabel metal1 2438 9486 2438 9486 0 ConfigBits\[7\]
rlabel metal2 8418 21692 8418 21692 0 ConfigBits\[80\]
rlabel metal2 9200 22406 9200 22406 0 ConfigBits\[81\]
rlabel metal1 11638 22474 11638 22474 0 ConfigBits\[82\]
rlabel metal2 12742 22950 12742 22950 0 ConfigBits\[83\]
rlabel metal1 7590 24344 7590 24344 0 ConfigBits\[84\]
rlabel metal1 8372 24242 8372 24242 0 ConfigBits\[85\]
rlabel metal1 12880 29070 12880 29070 0 ConfigBits\[86\]
rlabel via1 12189 29138 12189 29138 0 ConfigBits\[87\]
rlabel metal1 8372 30090 8372 30090 0 ConfigBits\[88\]
rlabel metal2 9430 31212 9430 31212 0 ConfigBits\[89\]
rlabel metal1 11546 18224 11546 18224 0 ConfigBits\[8\]
rlabel viali 12653 31858 12653 31858 0 ConfigBits\[90\]
rlabel metal2 13202 31841 13202 31841 0 ConfigBits\[91\]
rlabel metal1 7084 20978 7084 20978 0 ConfigBits\[92\]
rlabel metal1 7314 21862 7314 21862 0 ConfigBits\[93\]
rlabel metal1 12650 32232 12650 32232 0 ConfigBits\[94\]
rlabel metal1 13478 30770 13478 30770 0 ConfigBits\[95\]
rlabel metal1 8556 29070 8556 29070 0 ConfigBits\[96\]
rlabel metal2 8050 31969 8050 31969 0 ConfigBits\[97\]
rlabel metal1 11960 33830 11960 33830 0 ConfigBits\[98\]
rlabel metal2 12650 32436 12650 32436 0 ConfigBits\[99\]
rlabel metal1 6854 18768 6854 18768 0 ConfigBits\[9\]
rlabel metal1 13892 17306 13892 17306 0 E1BEG[0]
rlabel metal3 15717 18564 15717 18564 0 E1BEG[1]
rlabel metal3 15004 18836 15004 18836 0 E1BEG[2]
rlabel metal1 13386 18938 13386 18938 0 E1BEG[3]
rlabel metal3 14866 19380 14866 19380 0 E2BEG[0]
rlabel metal1 14950 17306 14950 17306 0 E2BEG[1]
rlabel metal3 14912 19924 14912 19924 0 E2BEG[2]
rlabel metal2 14398 19839 14398 19839 0 E2BEG[3]
rlabel metal3 14222 20468 14222 20468 0 E2BEG[4]
rlabel metal3 15533 20740 15533 20740 0 E2BEG[5]
rlabel metal3 15096 21012 15096 21012 0 E2BEG[6]
rlabel metal3 15073 21284 15073 21284 0 E2BEG[7]
rlabel metal3 15004 21556 15004 21556 0 E2BEGb[0]
rlabel metal1 14628 20570 14628 20570 0 E2BEGb[1]
rlabel metal3 14866 22100 14866 22100 0 E2BEGb[2]
rlabel metal1 12558 21624 12558 21624 0 E2BEGb[3]
rlabel metal2 14306 22423 14306 22423 0 E2BEGb[4]
rlabel metal3 15510 22916 15510 22916 0 E2BEGb[5]
rlabel metal1 14352 22746 14352 22746 0 E2BEGb[6]
rlabel metal3 15050 23460 15050 23460 0 E2BEGb[7]
rlabel metal3 15809 28084 15809 28084 0 E6BEG[0]
rlabel metal1 14260 32810 14260 32810 0 E6BEG[10]
rlabel metal3 15073 31076 15073 31076 0 E6BEG[11]
rlabel metal1 14766 32198 14766 32198 0 E6BEG[1]
rlabel metal1 14076 32334 14076 32334 0 E6BEG[2]
rlabel metal3 14981 28900 14981 28900 0 E6BEG[3]
rlabel metal3 14866 29172 14866 29172 0 E6BEG[4]
rlabel metal3 15533 29444 15533 29444 0 E6BEG[5]
rlabel metal3 15625 29716 15625 29716 0 E6BEG[6]
rlabel metal3 15050 29988 15050 29988 0 E6BEG[7]
rlabel metal1 13432 32198 13432 32198 0 E6BEG[8]
rlabel metal1 15088 34578 15088 34578 0 E6BEG[9]
rlabel metal3 15165 23732 15165 23732 0 EE4BEG[0]
rlabel metal2 11914 27421 11914 27421 0 EE4BEG[10]
rlabel metal3 15280 26724 15280 26724 0 EE4BEG[11]
rlabel metal3 15050 26996 15050 26996 0 EE4BEG[12]
rlabel metal3 15533 27268 15533 27268 0 EE4BEG[13]
rlabel metal3 15694 27540 15694 27540 0 EE4BEG[14]
rlabel metal3 14705 27812 14705 27812 0 EE4BEG[15]
rlabel metal3 15510 24004 15510 24004 0 EE4BEG[1]
rlabel metal2 12006 24735 12006 24735 0 EE4BEG[2]
rlabel metal3 15349 24548 15349 24548 0 EE4BEG[3]
rlabel metal2 11914 25245 11914 25245 0 EE4BEG[4]
rlabel metal3 15533 25092 15533 25092 0 EE4BEG[5]
rlabel metal3 15809 25364 15809 25364 0 EE4BEG[6]
rlabel metal3 15050 25636 15050 25636 0 EE4BEG[7]
rlabel metal3 15694 25908 15694 25908 0 EE4BEG[8]
rlabel metal3 15510 26180 15510 26180 0 EE4BEG[9]
rlabel metal3 452 15572 452 15572 0 FrameData[0]
rlabel metal3 452 23732 452 23732 0 FrameData[10]
rlabel metal3 452 24548 452 24548 0 FrameData[11]
rlabel metal3 452 25364 452 25364 0 FrameData[12]
rlabel metal3 820 26180 820 26180 0 FrameData[13]
rlabel metal3 452 26996 452 26996 0 FrameData[14]
rlabel metal3 452 27812 452 27812 0 FrameData[15]
rlabel metal3 452 28628 452 28628 0 FrameData[16]
rlabel metal3 452 29444 452 29444 0 FrameData[17]
rlabel metal3 774 30260 774 30260 0 FrameData[18]
rlabel metal3 452 31076 452 31076 0 FrameData[19]
rlabel metal3 475 16388 475 16388 0 FrameData[1]
rlabel metal3 452 31892 452 31892 0 FrameData[20]
rlabel metal3 452 32708 452 32708 0 FrameData[21]
rlabel metal3 452 33524 452 33524 0 FrameData[22]
rlabel metal3 452 34340 452 34340 0 FrameData[23]
rlabel metal3 452 35156 452 35156 0 FrameData[24]
rlabel metal3 452 35972 452 35972 0 FrameData[25]
rlabel metal3 452 36788 452 36788 0 FrameData[26]
rlabel metal3 452 37604 452 37604 0 FrameData[27]
rlabel metal3 475 38420 475 38420 0 FrameData[28]
rlabel metal3 452 39236 452 39236 0 FrameData[29]
rlabel metal3 452 17204 452 17204 0 FrameData[2]
rlabel metal3 452 40052 452 40052 0 FrameData[30]
rlabel metal3 452 40868 452 40868 0 FrameData[31]
rlabel metal3 452 18020 452 18020 0 FrameData[3]
rlabel metal3 820 18836 820 18836 0 FrameData[4]
rlabel metal3 452 19652 452 19652 0 FrameData[5]
rlabel metal3 452 20468 452 20468 0 FrameData[6]
rlabel metal3 452 21284 452 21284 0 FrameData[7]
rlabel metal3 452 22100 452 22100 0 FrameData[8]
rlabel metal3 452 22916 452 22916 0 FrameData[9]
rlabel metal3 15740 31348 15740 31348 0 FrameData_O[0]
rlabel metal3 14590 34068 14590 34068 0 FrameData_O[10]
rlabel metal3 15809 34340 15809 34340 0 FrameData_O[11]
rlabel metal3 14866 34612 14866 34612 0 FrameData_O[12]
rlabel metal3 15510 34884 15510 34884 0 FrameData_O[13]
rlabel metal3 15188 35156 15188 35156 0 FrameData_O[14]
rlabel metal3 15165 35428 15165 35428 0 FrameData_O[15]
rlabel metal3 15717 35700 15717 35700 0 FrameData_O[16]
rlabel metal3 15510 35972 15510 35972 0 FrameData_O[17]
rlabel metal3 14866 36244 14866 36244 0 FrameData_O[18]
rlabel metal3 15142 36516 15142 36516 0 FrameData_O[19]
rlabel metal1 14950 35462 14950 35462 0 FrameData_O[1]
rlabel metal3 14820 36788 14820 36788 0 FrameData_O[20]
rlabel metal3 15533 37060 15533 37060 0 FrameData_O[21]
rlabel metal3 14958 37332 14958 37332 0 FrameData_O[22]
rlabel metal3 15142 37604 15142 37604 0 FrameData_O[23]
rlabel metal3 14866 37876 14866 37876 0 FrameData_O[24]
rlabel metal3 15533 38148 15533 38148 0 FrameData_O[25]
rlabel metal3 15441 38420 15441 38420 0 FrameData_O[26]
rlabel metal3 15142 38692 15142 38692 0 FrameData_O[27]
rlabel metal3 14912 38964 14912 38964 0 FrameData_O[28]
rlabel metal3 15533 39236 15533 39236 0 FrameData_O[29]
rlabel metal3 15073 31892 15073 31892 0 FrameData_O[2]
rlabel metal3 15050 39508 15050 39508 0 FrameData_O[30]
rlabel metal3 14820 39780 14820 39780 0 FrameData_O[31]
rlabel metal3 15740 32164 15740 32164 0 FrameData_O[3]
rlabel metal2 12374 33473 12374 33473 0 FrameData_O[4]
rlabel metal3 15533 32708 15533 32708 0 FrameData_O[5]
rlabel metal3 14774 32980 14774 32980 0 FrameData_O[6]
rlabel metal3 14866 33252 14866 33252 0 FrameData_O[7]
rlabel metal3 15533 33524 15533 33524 0 FrameData_O[8]
rlabel metal3 15717 33796 15717 33796 0 FrameData_O[9]
rlabel metal1 11408 30090 11408 30090 0 FrameData_O_i\[0\]
rlabel metal1 12926 35156 12926 35156 0 FrameData_O_i\[10\]
rlabel metal1 11362 35598 11362 35598 0 FrameData_O_i\[11\]
rlabel metal2 10534 34340 10534 34340 0 FrameData_O_i\[12\]
rlabel metal1 12558 36652 12558 36652 0 FrameData_O_i\[13\]
rlabel metal2 10258 34952 10258 34952 0 FrameData_O_i\[14\]
rlabel metal2 10994 34884 10994 34884 0 FrameData_O_i\[15\]
rlabel metal1 12696 36346 12696 36346 0 FrameData_O_i\[16\]
rlabel metal1 11822 35666 11822 35666 0 FrameData_O_i\[17\]
rlabel metal1 9844 35258 9844 35258 0 FrameData_O_i\[18\]
rlabel metal1 8878 35802 8878 35802 0 FrameData_O_i\[19\]
rlabel metal1 10718 31858 10718 31858 0 FrameData_O_i\[1\]
rlabel metal1 13386 36312 13386 36312 0 FrameData_O_i\[20\]
rlabel metal1 11868 36346 11868 36346 0 FrameData_O_i\[21\]
rlabel metal1 12880 37230 12880 37230 0 FrameData_O_i\[22\]
rlabel metal1 12466 36856 12466 36856 0 FrameData_O_i\[23\]
rlabel metal1 13202 38896 13202 38896 0 FrameData_O_i\[24\]
rlabel metal1 12834 37876 12834 37876 0 FrameData_O_i\[25\]
rlabel metal2 10810 37638 10810 37638 0 FrameData_O_i\[26\]
rlabel metal2 12650 38148 12650 38148 0 FrameData_O_i\[27\]
rlabel metal2 12742 38726 12742 38726 0 FrameData_O_i\[28\]
rlabel metal1 13202 39372 13202 39372 0 FrameData_O_i\[29\]
rlabel metal1 10902 31790 10902 31790 0 FrameData_O_i\[2\]
rlabel metal1 9706 39440 9706 39440 0 FrameData_O_i\[30\]
rlabel metal1 10258 40052 10258 40052 0 FrameData_O_i\[31\]
rlabel metal1 11178 31790 11178 31790 0 FrameData_O_i\[3\]
rlabel metal1 14214 31994 14214 31994 0 FrameData_O_i\[4\]
rlabel metal1 12029 32878 12029 32878 0 FrameData_O_i\[5\]
rlabel metal2 8970 32436 8970 32436 0 FrameData_O_i\[6\]
rlabel metal1 10718 32912 10718 32912 0 FrameData_O_i\[7\]
rlabel metal1 11546 33082 11546 33082 0 FrameData_O_i\[8\]
rlabel metal2 10902 35343 10902 35343 0 FrameData_O_i\[9\]
rlabel metal2 1334 1010 1334 1010 0 FrameStrobe[0]
rlabel metal2 8694 704 8694 704 0 FrameStrobe[10]
rlabel metal2 9575 68 9575 68 0 FrameStrobe[11]
rlabel metal2 10166 704 10166 704 0 FrameStrobe[12]
rlabel metal2 10902 704 10902 704 0 FrameStrobe[13]
rlabel metal2 11638 704 11638 704 0 FrameStrobe[14]
rlabel metal2 12374 704 12374 704 0 FrameStrobe[15]
rlabel metal2 13110 143 13110 143 0 FrameStrobe[16]
rlabel metal2 13899 68 13899 68 0 FrameStrobe[17]
rlabel metal2 14582 704 14582 704 0 FrameStrobe[18]
rlabel metal2 15318 636 15318 636 0 FrameStrobe[19]
rlabel metal2 2070 704 2070 704 0 FrameStrobe[1]
rlabel metal2 2951 68 2951 68 0 FrameStrobe[2]
rlabel metal2 3687 68 3687 68 0 FrameStrobe[3]
rlabel metal2 4278 670 4278 670 0 FrameStrobe[4]
rlabel metal2 5113 68 5113 68 0 FrameStrobe[5]
rlabel metal2 5750 704 5750 704 0 FrameStrobe[6]
rlabel metal2 6486 704 6486 704 0 FrameStrobe[7]
rlabel metal2 7222 704 7222 704 0 FrameStrobe[8]
rlabel metal2 7958 143 7958 143 0 FrameStrobe[9]
rlabel metal2 1479 44948 1479 44948 0 FrameStrobe_O[0]
rlabel metal1 8924 43418 8924 43418 0 FrameStrobe_O[10]
rlabel metal2 9430 44176 9430 44176 0 FrameStrobe_O[11]
rlabel metal2 10442 44183 10442 44183 0 FrameStrobe_O[12]
rlabel metal2 10902 44176 10902 44176 0 FrameStrobe_O[13]
rlabel metal1 12098 43418 12098 43418 0 FrameStrobe_O[14]
rlabel metal2 12374 44176 12374 44176 0 FrameStrobe_O[15]
rlabel metal1 13202 43418 13202 43418 0 FrameStrobe_O[16]
rlabel metal2 13846 43632 13846 43632 0 FrameStrobe_O[17]
rlabel metal1 14214 42738 14214 42738 0 FrameStrobe_O[18]
rlabel metal1 14582 43418 14582 43418 0 FrameStrobe_O[19]
rlabel metal2 2346 44183 2346 44183 0 FrameStrobe_O[1]
rlabel metal2 2859 44948 2859 44948 0 FrameStrobe_O[2]
rlabel metal1 3772 43418 3772 43418 0 FrameStrobe_O[3]
rlabel metal2 4278 44176 4278 44176 0 FrameStrobe_O[4]
rlabel metal2 5290 44183 5290 44183 0 FrameStrobe_O[5]
rlabel metal2 5849 44948 5849 44948 0 FrameStrobe_O[6]
rlabel metal2 6631 44948 6631 44948 0 FrameStrobe_O[7]
rlabel metal2 7498 44183 7498 44183 0 FrameStrobe_O[8]
rlabel metal2 8103 44948 8103 44948 0 FrameStrobe_O[9]
rlabel metal1 1794 35258 1794 35258 0 FrameStrobe_O_i\[0\]
rlabel metal1 5405 42262 5405 42262 0 FrameStrobe_O_i\[10\]
rlabel metal1 9154 2074 9154 2074 0 FrameStrobe_O_i\[11\]
rlabel metal1 10120 2074 10120 2074 0 FrameStrobe_O_i\[12\]
rlabel metal3 11017 2652 11017 2652 0 FrameStrobe_O_i\[13\]
rlabel metal1 11776 2074 11776 2074 0 FrameStrobe_O_i\[14\]
rlabel via2 12466 42653 12466 42653 0 FrameStrobe_O_i\[15\]
rlabel metal1 14306 1802 14306 1802 0 FrameStrobe_O_i\[16\]
rlabel metal1 14582 1870 14582 1870 0 FrameStrobe_O_i\[17\]
rlabel metal2 13938 41797 13938 41797 0 FrameStrobe_O_i\[18\]
rlabel metal1 14858 1258 14858 1258 0 FrameStrobe_O_i\[19\]
rlabel metal1 2162 32538 2162 32538 0 FrameStrobe_O_i\[1\]
rlabel metal1 2990 26554 2990 26554 0 FrameStrobe_O_i\[2\]
rlabel metal2 3358 21597 3358 21597 0 FrameStrobe_O_i\[3\]
rlabel metal2 4094 42500 4094 42500 0 FrameStrobe_O_i\[4\]
rlabel metal1 5014 42330 5014 42330 0 FrameStrobe_O_i\[5\]
rlabel metal1 4922 42534 4922 42534 0 FrameStrobe_O_i\[6\]
rlabel metal1 5198 42738 5198 42738 0 FrameStrobe_O_i\[7\]
rlabel metal1 5497 2006 5497 2006 0 FrameStrobe_O_i\[8\]
rlabel metal1 1380 11594 1380 11594 0 FrameStrobe_O_i\[9\]
rlabel metal1 11270 7514 11270 7514 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out0
rlabel metal1 11132 8942 11132 8942 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out1
rlabel metal1 13386 9078 13386 9078 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out2
rlabel metal1 11730 9010 11730 9010 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out3
rlabel metal1 11546 6222 11546 6222 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out0
rlabel metal1 11546 6324 11546 6324 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out1
rlabel via1 12570 6290 12570 6290 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out2
rlabel via2 12466 6307 12466 6307 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out3
rlabel metal2 14122 18496 14122 18496 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN\[0\]
rlabel metal1 12190 18292 12190 18292 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN\[1\]
rlabel metal1 12006 18122 12006 18122 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_0_
rlabel metal1 11960 18190 11960 18190 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_1_
rlabel metal1 7590 18768 7590 18768 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN\[0\]
rlabel metal1 6900 19414 6900 19414 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN\[1\]
rlabel metal1 7314 18666 7314 18666 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_0_
rlabel metal1 7130 18836 7130 18836 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_1_
rlabel metal1 7406 19346 7406 19346 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN\[0\]
rlabel metal1 7498 20468 7498 20468 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN\[1\]
rlabel metal1 7406 19210 7406 19210 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_0_
rlabel via1 7407 19278 7407 19278 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_1_
rlabel metal1 10856 19346 10856 19346 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN\[0\]
rlabel metal1 11362 20468 11362 20468 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN\[1\]
rlabel metal1 11270 19210 11270 19210 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_0_
rlabel metal1 11776 19278 11776 19278 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_1_
rlabel metal1 6486 8500 6486 8500 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN\[0\]
rlabel metal2 6946 9078 6946 9078 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN\[1\]
rlabel metal1 6624 8602 6624 8602 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_0_
rlabel metal1 6716 9010 6716 9010 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_1_
rlabel metal1 6210 8432 6210 8432 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out0
rlabel metal1 7360 8466 7360 8466 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out1
rlabel metal1 7636 10234 7636 10234 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN\[0\]
rlabel metal1 7268 10030 7268 10030 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN\[1\]
rlabel metal1 5934 10574 5934 10574 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_0_
rlabel metal1 6210 10540 6210 10540 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_1_
rlabel metal1 8418 10030 8418 10030 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out0
rlabel metal1 7774 10064 7774 10064 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out1
rlabel metal1 3128 42602 3128 42602 0 UserCLK
rlabel metal1 3450 43384 3450 43384 0 UserCLKo
rlabel metal3 14820 5236 14820 5236 0 W1END[0]
rlabel metal3 15510 5508 15510 5508 0 W1END[1]
rlabel metal3 15441 5780 15441 5780 0 W1END[2]
rlabel metal3 15050 6052 15050 6052 0 W1END[3]
rlabel metal1 11132 7922 11132 7922 0 W2END[0]
rlabel metal3 15510 8772 15510 8772 0 W2END[1]
rlabel metal3 14337 9044 14337 9044 0 W2END[2]
rlabel metal3 14866 9316 14866 9316 0 W2END[3]
rlabel metal3 15096 9588 15096 9588 0 W2END[4]
rlabel metal3 15694 9860 15694 9860 0 W2END[5]
rlabel metal3 15510 10132 15510 10132 0 W2END[6]
rlabel metal3 15050 10404 15050 10404 0 W2END[7]
rlabel metal1 14214 6290 14214 6290 0 W2MID[0]
rlabel metal3 15510 6596 15510 6596 0 W2MID[1]
rlabel metal2 12374 5219 12374 5219 0 W2MID[2]
rlabel metal2 13662 4403 13662 4403 0 W2MID[3]
rlabel metal3 14820 7412 14820 7412 0 W2MID[4]
rlabel metal3 15510 7684 15510 7684 0 W2MID[5]
rlabel metal3 14636 7956 14636 7956 0 W2MID[6]
rlabel metal3 15096 8228 15096 8228 0 W2MID[7]
rlabel metal3 13946 15028 13946 15028 0 W6END[0]
rlabel metal2 11178 18003 11178 18003 0 W6END[10]
rlabel metal3 15073 18020 15073 18020 0 W6END[11]
rlabel metal3 15533 15300 15533 15300 0 W6END[1]
rlabel metal3 14590 15572 14590 15572 0 W6END[2]
rlabel metal3 15786 15844 15786 15844 0 W6END[3]
rlabel metal3 15050 16116 15050 16116 0 W6END[4]
rlabel metal3 15533 16388 15533 16388 0 W6END[5]
rlabel metal3 15096 16660 15096 16660 0 W6END[6]
rlabel metal3 15234 16932 15234 16932 0 W6END[7]
rlabel metal3 13808 17204 13808 17204 0 W6END[8]
rlabel metal3 15556 17476 15556 17476 0 W6END[9]
rlabel metal2 11086 10897 11086 10897 0 WW4END[0]
rlabel metal3 15050 13396 15050 13396 0 WW4END[10]
rlabel metal3 15280 13668 15280 13668 0 WW4END[11]
rlabel metal3 14820 13940 14820 13940 0 WW4END[12]
rlabel metal3 15809 14212 15809 14212 0 WW4END[13]
rlabel metal3 15694 14484 15694 14484 0 WW4END[14]
rlabel metal3 15096 14756 15096 14756 0 WW4END[15]
rlabel metal3 15533 10948 15533 10948 0 WW4END[1]
rlabel metal1 11546 11118 11546 11118 0 WW4END[2]
rlabel metal3 15280 11492 15280 11492 0 WW4END[3]
rlabel metal3 15050 11764 15050 11764 0 WW4END[4]
rlabel metal3 15510 12036 15510 12036 0 WW4END[5]
rlabel metal2 11822 12563 11822 12563 0 WW4END[6]
rlabel metal3 14912 12580 14912 12580 0 WW4END[7]
rlabel metal1 13570 12274 13570 12274 0 WW4END[8]
rlabel metal3 15556 13124 15556 13124 0 WW4END[9]
rlabel metal1 4544 18258 4544 18258 0 net1
rlabel metal2 2024 16560 2024 16560 0 net10
rlabel metal1 12535 21454 12535 21454 0 net100
rlabel via2 12006 31773 12006 31773 0 net101
rlabel metal1 12512 12614 12512 12614 0 net102
rlabel metal1 1564 10778 1564 10778 0 net103
rlabel metal2 2438 10642 2438 10642 0 net104
rlabel metal1 1748 12138 1748 12138 0 net105
rlabel metal1 1748 13294 1748 13294 0 net106
rlabel metal1 1748 13974 1748 13974 0 net107
rlabel metal1 1656 15062 1656 15062 0 net108
rlabel metal1 1932 5610 1932 5610 0 net109
rlabel metal1 1747 16558 1747 16558 0 net11
rlabel metal1 1840 5270 1840 5270 0 net110
rlabel metal1 2162 6664 2162 6664 0 net111
rlabel metal1 1978 6970 1978 6970 0 net112
rlabel metal1 1518 8568 1518 8568 0 net113
rlabel metal2 2806 9826 2806 9826 0 net114
rlabel metal1 13478 17170 13478 17170 0 net115
rlabel metal1 7130 17612 7130 17612 0 net116
rlabel metal1 10718 19346 10718 19346 0 net117
rlabel metal1 12190 18768 12190 18768 0 net118
rlabel metal1 9154 17306 9154 17306 0 net119
rlabel metal1 5658 13770 5658 13770 0 net12
rlabel metal1 12971 17238 12971 17238 0 net120
rlabel metal2 10442 16609 10442 16609 0 net121
rlabel metal2 14490 18870 14490 18870 0 net122
rlabel metal1 12236 14586 12236 14586 0 net123
rlabel metal1 13156 13498 13156 13498 0 net124
rlabel metal1 10856 20026 10856 20026 0 net125
rlabel metal1 13846 16694 13846 16694 0 net126
rlabel metal1 12834 20876 12834 20876 0 net127
rlabel metal2 11638 21182 11638 21182 0 net128
rlabel metal2 13570 22559 13570 22559 0 net129
rlabel metal1 1426 31110 1426 31110 0 net13
rlabel metal1 13892 20026 13892 20026 0 net130
rlabel metal2 14352 20332 14352 20332 0 net131
rlabel metal1 15042 11866 15042 11866 0 net132
rlabel metal2 12466 15402 12466 15402 0 net133
rlabel metal2 12190 22899 12190 22899 0 net134
rlabel metal1 11592 29818 11592 29818 0 net135
rlabel metal2 13018 32640 13018 32640 0 net136
rlabel metal1 13294 31382 13294 31382 0 net137
rlabel metal2 14122 32071 14122 32071 0 net138
rlabel metal1 14260 31926 14260 31926 0 net139
rlabel metal1 1656 17306 1656 17306 0 net14
rlabel metal1 10672 30226 10672 30226 0 net140
rlabel metal1 9062 24038 9062 24038 0 net141
rlabel metal1 11316 29206 11316 29206 0 net142
rlabel metal1 10534 30294 10534 30294 0 net143
rlabel metal2 11546 31841 11546 31841 0 net144
rlabel metal2 13018 32351 13018 32351 0 net145
rlabel metal2 14030 33388 14030 33388 0 net146
rlabel metal1 13110 24378 13110 24378 0 net147
rlabel metal2 13386 27710 13386 27710 0 net148
rlabel metal1 13616 26554 13616 26554 0 net149
rlabel viali 1693 8912 1693 8912 0 net15
rlabel metal1 11040 27438 11040 27438 0 net150
rlabel metal2 10534 29444 10534 29444 0 net151
rlabel metal2 13846 21556 13846 21556 0 net152
rlabel metal1 14766 33490 14766 33490 0 net153
rlabel metal1 14398 23766 14398 23766 0 net154
rlabel metal2 8234 24480 8234 24480 0 net155
rlabel metal2 13754 27880 13754 27880 0 net156
rlabel metal2 5198 17204 5198 17204 0 net157
rlabel via2 14490 12699 14490 12699 0 net158
rlabel metal2 14582 17476 14582 17476 0 net159
rlabel metal1 1747 9554 1747 9554 0 net16
rlabel metal1 14858 15402 14858 15402 0 net160
rlabel metal1 14306 26010 14306 26010 0 net161
rlabel metal1 8740 29546 8740 29546 0 net162
rlabel metal1 12719 32878 12719 32878 0 net163
rlabel viali 13018 35052 13018 35052 0 net164
rlabel metal2 13202 35836 13202 35836 0 net165
rlabel metal2 13570 35190 13570 35190 0 net166
rlabel metal2 12466 36142 12466 36142 0 net167
rlabel metal1 13018 35768 13018 35768 0 net168
rlabel metal2 12834 35411 12834 35411 0 net169
rlabel via2 13110 37213 13110 37213 0 net17
rlabel metal1 12926 36890 12926 36890 0 net170
rlabel metal1 11546 35768 11546 35768 0 net171
rlabel metal1 12466 36720 12466 36720 0 net172
rlabel metal1 13478 37196 13478 37196 0 net173
rlabel metal2 13662 35343 13662 35343 0 net174
rlabel metal1 13386 37434 13386 37434 0 net175
rlabel metal1 14122 37774 14122 37774 0 net176
rlabel metal2 12650 37604 12650 37604 0 net177
rlabel metal1 14214 38284 14214 38284 0 net178
rlabel metal1 13754 38318 13754 38318 0 net179
rlabel metal2 12834 5168 12834 5168 0 net18
rlabel metal1 13018 37638 13018 37638 0 net180
rlabel metal1 12742 37944 12742 37944 0 net181
rlabel metal1 12880 38454 12880 38454 0 net182
rlabel metal1 13156 39066 13156 39066 0 net183
rlabel metal1 13202 39610 13202 39610 0 net184
rlabel metal2 10810 32776 10810 32776 0 net185
rlabel metal2 13938 39780 13938 39780 0 net186
rlabel metal2 13570 40290 13570 40290 0 net187
rlabel metal1 11730 31994 11730 31994 0 net188
rlabel metal1 13294 33082 13294 33082 0 net189
rlabel metal2 12558 36193 12558 36193 0 net19
rlabel metal1 11776 32742 11776 32742 0 net190
rlabel metal2 13294 36465 13294 36465 0 net191
rlabel via2 13570 34595 13570 34595 0 net192
rlabel metal1 12995 34986 12995 34986 0 net193
rlabel metal1 11316 34646 11316 34646 0 net194
rlabel metal1 1656 43282 1656 43282 0 net195
rlabel metal1 8786 42874 8786 42874 0 net196
rlabel metal2 9246 43078 9246 43078 0 net197
rlabel metal2 10258 43078 10258 43078 0 net198
rlabel metal1 11224 42874 11224 42874 0 net199
rlabel metal2 3910 7922 3910 7922 0 net2
rlabel metal2 13478 37485 13478 37485 0 net20
rlabel metal1 11822 42806 11822 42806 0 net200
rlabel metal1 12420 42874 12420 42874 0 net201
rlabel metal1 12926 42874 12926 42874 0 net202
rlabel metal2 14122 42670 14122 42670 0 net203
rlabel metal1 13662 42330 13662 42330 0 net204
rlabel metal1 13938 42534 13938 42534 0 net205
rlabel metal1 2116 42330 2116 42330 0 net206
rlabel metal1 2944 43282 2944 43282 0 net207
rlabel metal1 3588 42874 3588 42874 0 net208
rlabel metal1 4324 42874 4324 42874 0 net209
rlabel viali 6477 17616 6477 17616 0 net21
rlabel metal1 5014 42874 5014 42874 0 net210
rlabel metal1 5750 42874 5750 42874 0 net211
rlabel metal1 6532 42874 6532 42874 0 net212
rlabel metal1 7222 42874 7222 42874 0 net213
rlabel metal1 8004 42874 8004 42874 0 net214
rlabel metal1 3082 42874 3082 42874 0 net215
rlabel metal1 8303 8398 8303 8398 0 net216
rlabel metal1 8165 10574 8165 10574 0 net217
rlabel metal2 8326 8976 8326 8976 0 net218
rlabel metal1 7222 10574 7222 10574 0 net219
rlabel metal1 7957 16558 7957 16558 0 net22
rlabel metal1 12880 38318 12880 38318 0 net23
rlabel metal2 1610 39168 1610 39168 0 net24
rlabel metal1 6715 24786 6715 24786 0 net25
rlabel metal1 7067 16082 7067 16082 0 net26
rlabel via1 9245 15470 9245 15470 0 net27
rlabel metal1 1702 18088 1702 18088 0 net28
rlabel metal3 10235 18700 10235 18700 0 net29
rlabel metal2 8418 17255 8418 17255 0 net3
rlabel metal2 5612 20740 5612 20740 0 net30
rlabel metal1 7313 30226 7313 30226 0 net31
rlabel metal1 8463 20434 8463 20434 0 net32
rlabel metal1 1656 22746 1656 22746 0 net33
rlabel metal2 14030 35122 14030 35122 0 net34
rlabel metal1 2254 1836 2254 1836 0 net35
rlabel metal1 8786 1530 8786 1530 0 net36
rlabel metal1 9430 1530 9430 1530 0 net37
rlabel metal1 10212 1530 10212 1530 0 net38
rlabel metal1 10948 1530 10948 1530 0 net39
rlabel viali 12434 21968 12434 21968 0 net4
rlabel metal1 11684 1530 11684 1530 0 net40
rlabel metal1 12420 1530 12420 1530 0 net41
rlabel metal1 13248 1530 13248 1530 0 net42
rlabel metal2 13754 1734 13754 1734 0 net43
rlabel metal2 13478 1768 13478 1768 0 net44
rlabel metal1 13708 1258 13708 1258 0 net45
rlabel metal1 7774 1394 7774 1394 0 net46
rlabel metal1 7452 1870 7452 1870 0 net47
rlabel metal1 1518 6290 1518 6290 0 net48
rlabel via2 4646 1309 4646 1309 0 net49
rlabel metal2 12834 21284 12834 21284 0 net5
rlabel via2 5382 1309 5382 1309 0 net50
rlabel metal1 5796 1530 5796 1530 0 net51
rlabel metal1 6532 1530 6532 1530 0 net52
rlabel metal1 7268 1530 7268 1530 0 net53
rlabel metal1 8004 1530 8004 1530 0 net54
rlabel metal2 14306 11152 14306 11152 0 net55
rlabel metal2 2484 16560 2484 16560 0 net56
rlabel metal1 7452 18734 7452 18734 0 net57
rlabel metal2 13570 28492 13570 28492 0 net58
rlabel metal1 7222 9010 7222 9010 0 net59
rlabel metal1 10057 32402 10057 32402 0 net6
rlabel metal2 11638 9486 11638 9486 0 net60
rlabel metal2 7866 9180 7866 9180 0 net61
rlabel metal1 7590 8364 7590 8364 0 net62
rlabel metal2 7406 9010 7406 9010 0 net63
rlabel metal1 6808 10574 6808 10574 0 net64
rlabel metal2 13478 9299 13478 9299 0 net65
rlabel metal1 14950 21930 14950 21930 0 net66
rlabel metal1 12098 16592 12098 16592 0 net67
rlabel via2 13662 6715 13662 6715 0 net68
rlabel metal1 13202 5644 13202 5644 0 net69
rlabel metal1 10073 25874 10073 25874 0 net7
rlabel metal1 10672 14450 10672 14450 0 net70
rlabel metal1 13754 9078 13754 9078 0 net71
rlabel metal2 13846 8160 13846 8160 0 net72
rlabel metal1 13478 7446 13478 7446 0 net73
rlabel metal2 13892 8364 13892 8364 0 net74
rlabel metal1 10994 24106 10994 24106 0 net75
rlabel via1 13674 23630 13674 23630 0 net76
rlabel metal1 11178 17850 11178 17850 0 net77
rlabel metal1 11500 15606 11500 15606 0 net78
rlabel metal1 11546 29036 11546 29036 0 net79
rlabel metal1 9614 33966 9614 33966 0 net8
rlabel metal1 13386 14280 13386 14280 0 net80
rlabel metal2 13248 30124 13248 30124 0 net81
rlabel metal1 6624 15062 6624 15062 0 net82
rlabel metal1 10626 22066 10626 22066 0 net83
rlabel metal1 13018 21454 13018 21454 0 net84
rlabel metal1 11730 17782 11730 17782 0 net85
rlabel via2 13846 17867 13846 17867 0 net86
rlabel metal2 11960 18700 11960 18700 0 net87
rlabel metal2 15824 23868 15824 23868 0 net88
rlabel metal1 13202 13192 13202 13192 0 net89
rlabel metal2 1472 21420 1472 21420 0 net9
rlabel via1 13674 18190 13674 18190 0 net90
rlabel metal1 6440 20910 6440 20910 0 net91
rlabel metal1 14490 16184 14490 16184 0 net92
rlabel metal1 15962 20740 15962 20740 0 net93
rlabel metal2 8970 20383 8970 20383 0 net94
rlabel metal2 13938 18700 13938 18700 0 net95
rlabel metal1 13340 11254 13340 11254 0 net96
rlabel metal1 11730 19890 11730 19890 0 net97
rlabel metal1 7222 14994 7222 14994 0 net98
rlabel metal2 9798 21879 9798 21879 0 net99
<< properties >>
string FIXED_BBOX 0 0 16000 45000
<< end >>
