* NGSPICE file created from RegFile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxbp_1 abstract view
.subckt sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

.subckt RegFile E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2] E1END[3]
+ E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0]
+ E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7] E2END[0] E2END[1]
+ E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2]
+ E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1]
+ E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] E6END[0]
+ E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5] E6END[6] E6END[7]
+ E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13] EE4BEG[14]
+ EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6] EE4BEG[7]
+ EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13] EE4END[14]
+ EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6] EE4END[7]
+ EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S1END[0]
+ S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5]
+ S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6]
+ S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7]
+ S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4BEG[0]
+ S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3]
+ S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0] W1BEG[1] W1BEG[2]
+ W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1] W2BEG[2] W2BEG[3]
+ W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2] W2BEGb[3] W2BEGb[4]
+ W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5]
+ W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6]
+ W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5]
+ W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11] W6END[1] W6END[2]
+ W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9] WW4BEG[0] WW4BEG[10]
+ WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1] WW4BEG[2] WW4BEG[3]
+ WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9] WW4END[0] WW4END[10]
+ WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1] WW4END[2] WW4END[3]
+ WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
XFILLER_0_76_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XW6END_inbuf_0__0_ net230 VGND VGND VPWR VPWR W6BEG_i\[0\] sky130_fd_sc_hd__clkbuf_2
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame1_bit9 net80 net92 VGND VGND VPWR VPWR ConfigBits\[359\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame11_bit5 net76 net83 VGND VGND VPWR VPWR ConfigBits\[35\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame7_bit18 net58 net98 VGND VGND VPWR VPWR ConfigBits\[176\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame0_bit20 net61 net81 VGND VGND VPWR VPWR ConfigBits\[402\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame0_bit31 net73 net81 VGND VGND VPWR VPWR ConfigBits\[413\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3/X ConfigBits\[112\]
+ ConfigBits\[113\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame7_bit29 net70 net98 VGND VGND VPWR VPWR ConfigBits\[187\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3/X ConfigBits\[332\]
+ ConfigBits\[333\] VGND VGND VPWR VPWR JS2BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XWW4END_inbuf_10__0_ net243 VGND VGND VPWR VPWR WW4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput401 net401 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1431_ net205 Inst_RegFile_32x4/_0083_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1431_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput434 net434 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput412 net412 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput423 net423 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1362_ net205 Inst_RegFile_32x4/_0022_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1362_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1293_ Inst_RegFile_32x4__1455_/Q Inst_RegFile_32x4/_0598_ Inst_RegFile_32x4/_0632_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0636_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix__01_ JE2BEG\[1\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__buf_1
Xoutput489 net489 VGND VGND VPWR VPWR W6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput445 net445 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput456 net456 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput467 net467 VGND VGND VPWR VPWR W2BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput478 net478 VGND VGND VPWR VPWR W2BEGb[7] sky130_fd_sc_hd__clkbuf_4
XN4BEG_outbuf_11__0_ N4BEG_i\[11\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame3_bit24 net65 net94 VGND VGND VPWR VPWR ConfigBits\[310\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit13 net53 net94 VGND VGND VPWR VPWR ConfigBits\[299\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4END_inbuf_9__0_ net177 VGND VGND VPWR VPWR S4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0931_ Inst_RegFile_32x4/_0385_ VGND VGND VPWR VPWR BD1 sky130_fd_sc_hd__buf_12
XFILLER_0_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0793_ Inst_RegFile_32x4__1407_/Q Inst_RegFile_32x4__1383_/Q Inst_RegFile_32x4/_0137_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0862_ Inst_RegFile_32x4/_0302_ Inst_RegFile_32x4/_0318_ Inst_RegFile_32x4/_0319_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0320_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput275 net275 VGND VGND VPWR VPWR E6BEG[10] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1414_ net205 Inst_RegFile_32x4/_0066_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1414_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput286 net286 VGND VGND VPWR VPWR EE4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput264 net264 VGND VGND VPWR VPWR E2BEG[6] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1345_ net205 Inst_RegFile_32x4/_0005_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1345_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput297 net297 VGND VGND VPWR VPWR EE4BEG[5] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1276_ Inst_RegFile_32x4/_0453_ Inst_RegFile_32x4/_0454_ Inst_RegFile_32x4/_0452_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0626_ sky130_fd_sc_hd__or3b_4
XFILLER_0_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG0 net112 net41 net164 net217
+ ConfigBits\[238\] ConfigBits\[239\] VGND VGND VPWR VPWR J2END_EF_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame7_bit4 net75 net98 VGND VGND VPWR VPWR ConfigBits\[162\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit17 net57 net97 VGND VGND VPWR VPWR ConfigBits\[207\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame6_bit28 net69 net97 VGND VGND VPWR VPWR ConfigBits\[218\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1130_ Inst_RegFile_32x4__1380_/Q Inst_RegFile_32x4/_0524_ Inst_RegFile_32x4/_0539_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1061_ Inst_RegFile_32x4/_0497_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0013_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0914_ Inst_RegFile_32x4/_0313_ Inst_RegFile_32x4/_0369_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0370_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0845_ Inst_RegFile_32x4/_0291_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0303_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame2_bit23 net64 net93 VGND VGND VPWR VPWR ConfigBits\[341\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0776_ Inst_RegFile_32x4__1450_/Q Inst_RegFile_32x4__1474_/Q Inst_RegFile_32x4/_0156_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0240_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame2_bit12 net52 net93 VGND VGND VPWR VPWR ConfigBits\[330\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1259_ Inst_RegFile_32x4__1440_/Q Inst_RegFile_32x4/_0591_ Inst_RegFile_32x4/_0616_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1328_ Inst_RegFile_32x4/_0655_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0122_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_my_mux2_inst__1_/A1 ConfigBits\[135\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_inbuf_20__0_ net61 VGND VGND VPWR VPWR FrameData_O_i\[20\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1113_ Inst_RegFile_32x4/_0529_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0033_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame5_bit27 net68 net96 VGND VGND VPWR VPWR ConfigBits\[249\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame5_bit16 net56 net96 VGND VGND VPWR VPWR ConfigBits\[238\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1044_ Inst_RegFile_32x4/_0483_ Inst_RegFile_32x4/_0485_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0486_ sky130_fd_sc_hd__nor2_2
Xdata_inbuf_11__0_ net51 VGND VGND VPWR VPWR FrameData_O_i\[11\] sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0828_ Inst_RegFile_32x4/_0287_ VGND VGND VPWR VPWR AD2 sky130_fd_sc_hd__buf_12
XInst_RegFile_ConfigMem_Inst_frame4_bit7 net78 net95 VGND VGND VPWR VPWR ConfigBits\[261\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0 net107
+ net129 net1 net7 ConfigBits\[258\] ConfigBits\[259\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0759_ Inst_RegFile_32x4__1358_/Q Inst_RegFile_32x4__1446_/Q Inst_RegFile_32x4/_0131_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_5 JN2BEG\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame1_bit22 net63 net92 VGND VGND VPWR VPWR ConfigBits\[372\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame1_bit11 net51 net92 VGND VGND VPWR VPWR ConfigBits\[361\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_S4BEG3 net158 net173 net226 AD3 ConfigBits\[72\]
+ ConfigBits\[73\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__mux4_1
XFILLER_0_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1027_ Inst_RegFile_32x4/_0472_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0473_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput197 SS4END[2] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_2
Xinput175 S4END[11] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
Xinput186 S4END[7] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xinput164 S2END[7] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_2
Xinput153 S1END[0] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
Xinput131 N4END[4] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
Xinput120 N2MID[7] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_4
Xinput142 NN4END[14] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_14__0_ FrameStrobe_O_i\[14\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3/X ConfigBits\[280\]
+ ConfigBits\[281\] VGND VGND VPWR VPWR JN2BEG\[6\] sky130_fd_sc_hd__mux4_2
XFILLER_0_66_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame4_bit26 net67 net95 VGND VGND VPWR VPWR ConfigBits\[280\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_9__0_ FrameData_O_i\[9\] VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame4_bit15 net55 net95 VGND VGND VPWR VPWR ConfigBits\[269\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame11_bit6 net77 net83 VGND VGND VPWR VPWR ConfigBits\[36\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XWW4END_inbuf_5__0_ net253 VGND VGND VPWR VPWR WW4BEG_i\[5\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst0 net103
+ net3 net155 AD1 ConfigBits\[38\] ConfigBits\[39\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame0_bit21 net62 net81 VGND VGND VPWR VPWR ConfigBits\[403\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame0_bit10 net50 net81 VGND VGND VPWR VPWR ConfigBits\[392\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame7_bit19 net59 net98 VGND VGND VPWR VPWR ConfigBits\[177\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput402 net402 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1292_ Inst_RegFile_32x4/_0635_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0106_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1430_ net205 Inst_RegFile_32x4/_0082_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1430_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1361_ net205 Inst_RegFile_32x4/_0021_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1361_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput446 net446 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput457 net457 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput435 net435 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput413 net413 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput424 net424 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput468 net468 VGND VGND VPWR VPWR W2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput479 net479 VGND VGND VPWR VPWR W6BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix__00_ JE2BEG\[0\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame3_bit25 net66 net94 VGND VGND VPWR VPWR ConfigBits\[311\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame3_bit14 net54 net94 VGND VGND VPWR VPWR ConfigBits\[300\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0930_ Inst_RegFile_32x4__1389_/D Inst_RegFile_32x4__1389_/Q ConfigBits\[1\]
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0385_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0861_ B_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0319_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0792_ Inst_RegFile_32x4/_0182_ Inst_RegFile_32x4/_0254_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0255_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1413_ net205 Inst_RegFile_32x4/_0065_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1413_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput276 net276 VGND VGND VPWR VPWR E6BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput287 net287 VGND VGND VPWR VPWR EE4BEG[10] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1275_ Inst_RegFile_32x4/_0625_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0099_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput298 net298 VGND VGND VPWR VPWR EE4BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput265 net265 VGND VGND VPWR VPWR E2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput254 net254 VGND VGND VPWR VPWR E1BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1344_ net205 Inst_RegFile_32x4/_0004_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1344_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG1 net108 net8 net160 net245
+ ConfigBits\[240\] ConfigBits\[241\] VGND VGND VPWR VPWR J2END_EF_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame7_bit5 net76 net98 VGND VGND VPWR VPWR ConfigBits\[163\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame6_bit29 net70 net97 VGND VGND VPWR VPWR ConfigBits\[219\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit18 net58 net97 VGND VGND VPWR VPWR ConfigBits\[208\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_inbuf_11__0_ net83 VGND VGND VPWR VPWR FrameStrobe_O_i\[11\] sky130_fd_sc_hd__clkbuf_1
XE6END_inbuf_5__0_ net30 VGND VGND VPWR VPWR E6BEG_i\[5\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1060_ Inst_RegFile_32x4__1353_/Q Inst_RegFile_32x4/_0496_ Inst_RegFile_32x4/_0494_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0913_ Inst_RegFile_32x4__1457_/Q Inst_RegFile_32x4__1453_/Q Inst_RegFile_32x4/_0326_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0844_ Inst_RegFile_32x4/_0289_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0302_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_70_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame2_bit24 net65 net93 VGND VGND VPWR VPWR ConfigBits\[342\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0775_ Inst_RegFile_32x4/_0152_ Inst_RegFile_32x4/_0238_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0239_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame2_bit13 net53 net93 VGND VGND VPWR VPWR ConfigBits\[331\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1258_ Inst_RegFile_32x4/_0474_ Inst_RegFile_32x4/_0600_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0616_ sky130_fd_sc_hd__and2_2
XInst_RegFile_32x4__1189_ Inst_RegFile_32x4/_0462_ Inst_RegFile_32x4__1413_/Q Inst_RegFile_32x4/_0572_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0574_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1327_ Inst_RegFile_32x4/_0479_ Inst_RegFile_32x4__1470_/Q Inst_RegFile_32x4/_0652_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0655_ sky130_fd_sc_hd__mux2_1
XSS4END_inbuf_7__0_ net191 VGND VGND VPWR VPWR SS4BEG_i\[7\] sky130_fd_sc_hd__buf_2
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame5_bit17 net57 net96 VGND VGND VPWR VPWR ConfigBits\[239\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1112_ Inst_RegFile_32x4__1373_/Q Inst_RegFile_32x4/_0528_ Inst_RegFile_32x4/_0526_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0529_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1043_ Inst_RegFile_32x4/_0456_ Inst_RegFile_32x4/_0484_ Inst_RegFile_32x4/_0457_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0485_ sky130_fd_sc_hd__nand3_4
Xstrobe_outbuf_9__0_ FrameStrobe_O_i\[9\] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame5_bit28 net69 net96 VGND VGND VPWR VPWR ConfigBits\[250\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1 net40
+ net21 net159 net212 ConfigBits\[258\] ConfigBits\[259\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame4_bit8 net79 net95 VGND VGND VPWR VPWR ConfigBits\[262\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0827_ Inst_RegFile_32x4__1386_/D Inst_RegFile_32x4__1386_/Q ConfigBits\[0\]
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0287_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0758_ Inst_RegFile_32x4/_0222_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1385_/D
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0689_ Inst_RegFile_32x4/_0152_ Inst_RegFile_32x4/_0154_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0155_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XEE4END_inbuf_6__0_ net34 VGND VGND VPWR VPWR EE4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_3__0_ net74 VGND VGND VPWR VPWR FrameData_O_i\[3\] sky130_fd_sc_hd__buf_1
XFILLER_0_53_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 JW2BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame1_bit23 net64 net92 VGND VGND VPWR VPWR ConfigBits\[373\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame1_bit12 net52 net92 VGND VGND VPWR VPWR ConfigBits\[362\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XWW4BEG_outbuf_7__0_ WW4BEG_i\[7\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0 net103
+ net109 net121 net9 ConfigBits\[298\] ConfigBits\[299\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1026_ W_ADR1 W_ADR0 W_en VGND VGND VPWR VPWR Inst_RegFile_32x4/_0472_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput110 N2END[5] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_2
Xinput198 SS4END[3] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_2
Xinput176 S4END[12] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xinput187 S4END[8] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
Xinput165 S2MID[0] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_2
Xinput154 S1END[1] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_4
Xinput132 N4END[5] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
Xinput121 N4END[0] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
Xinput143 NN4END[15] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame4_bit27 net68 net95 VGND VGND VPWR VPWR ConfigBits\[281\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame4_bit16 net56 net95 VGND VGND VPWR VPWR ConfigBits\[270\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4END_inbuf_9__0_ net125 VGND VGND VPWR VPWR N4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame11_bit7 net78 net83 VGND VGND VPWR VPWR ConfigBits\[37\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1009_ Inst_RegFile_32x4/_0455_ Inst_RegFile_32x4/_0458_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0459_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst1 BD1 J2MID_ABb_BEG\[1\]
+ J2MID_CDb_BEG\[1\] J2END_GH_BEG\[0\] ConfigBits\[38\] ConfigBits\[39\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame0_bit22 net63 net81 VGND VGND VPWR VPWR ConfigBits\[404\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame0_bit11 net51 net81 VGND VGND VPWR VPWR ConfigBits\[393\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst0 net101
+ net1 net206 AD3 ConfigBits\[24\] ConfigBits\[25\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XN4BEG_outbuf_1__0_ N4BEG_i\[1\] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame0_bit0 net49 net81 VGND VGND VPWR VPWR ConfigBits\[382\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput458 net458 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_2
Xoutput403 net403 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1291_ Inst_RegFile_32x4__1454_/Q Inst_RegFile_32x4/_0596_ Inst_RegFile_32x4/_0632_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0635_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0 net137
+ net4 net189 net209 ConfigBits\[50\] ConfigBits\[51\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1360_ net205 Inst_RegFile_32x4/_0020_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1360_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput447 net447 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput436 net436 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput414 net414 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput425 net425 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput469 net469 VGND VGND VPWR VPWR W2BEG[6] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG0 net119 net19 net171
+ JN2BEG\[6\] ConfigBits\[182\] ConfigBits\[183\] VGND VGND VPWR VPWR J2MID_GHa_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XSS4BEG_outbuf_0__0_ SS4BEG_i\[0\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame3_bit26 net67 net94 VGND VGND VPWR VPWR ConfigBits\[312\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit15 net55 net94 VGND VGND VPWR VPWR ConfigBits\[301\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix__59_ net221 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0 net103
+ net111 net3 net11 ConfigBits\[370\] ConfigBits\[371\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0791_ Inst_RegFile_32x4__1359_/Q Inst_RegFile_32x4__1447_/Q Inst_RegFile_32x4/_0131_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0254_ sky130_fd_sc_hd__mux2_1
XW6BEG_outbuf_1__0_ W6BEG_i\[1\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0860_ Inst_RegFile_32x4__1352_/Q Inst_RegFile_32x4__1348_/Q Inst_RegFile_32x4/_0317_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1412_ net205 Inst_RegFile_32x4/_0064_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1412_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput277 net277 VGND VGND VPWR VPWR E6BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput288 net288 VGND VGND VPWR VPWR EE4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput299 net299 VGND VGND VPWR VPWR EE4BEG[7] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1274_ Inst_RegFile_32x4__1447_/Q Inst_RegFile_32x4/_0598_ Inst_RegFile_32x4/_0621_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0625_ sky130_fd_sc_hd__mux2_1
Xoutput266 net266 VGND VGND VPWR VPWR E2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput255 net255 VGND VGND VPWR VPWR E1BEG[1] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1343_ net205 Inst_RegFile_32x4/_0003_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1343_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG2 net110 net10 net196 net215
+ ConfigBits\[242\] ConfigBits\[243\] VGND VGND VPWR VPWR J2END_EF_BEG\[2\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame7_bit6 net77 net98 VGND VGND VPWR VPWR ConfigBits\[164\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0989_ Inst_RegFile_32x4/_0434_ Inst_RegFile_32x4/_0436_ Inst_RegFile_32x4/_0438_
+ Inst_RegFile_32x4/_0440_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0441_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame6_bit19 net59 net97 VGND VGND VPWR VPWR ConfigBits\[209\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_30__0_ FrameData_O_i\[30\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0774_ Inst_RegFile_32x4__1458_/Q Inst_RegFile_32x4__1454_/Q Inst_RegFile_32x4/_0153_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0843_ Inst_RegFile_32x4/_0296_ Inst_RegFile_32x4/_0299_ Inst_RegFile_32x4/_0300_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0301_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0912_ Inst_RegFile_32x4/_0364_ Inst_RegFile_32x4/_0366_ Inst_RegFile_32x4/_0367_
+ Inst_RegFile_32x4/_0310_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0368_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame2_bit25 net66 net93 VGND VGND VPWR VPWR ConfigBits\[343\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame2_bit14 net54 net93 VGND VGND VPWR VPWR ConfigBits\[332\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1326_ Inst_RegFile_32x4/_0654_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0121_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_21__0_ FrameData_O_i\[21\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__1257_ Inst_RegFile_32x4/_0615_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0091_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1188_ Inst_RegFile_32x4/_0573_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0064_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0 net102
+ net110 net2 net10 ConfigBits\[334\] ConfigBits\[335\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_12__0_ FrameData_O_i\[12\] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XS4BEG_outbuf_1__0_ S4BEG_i\[1\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame5_bit18 net58 net96 VGND VGND VPWR VPWR ConfigBits\[240\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame5_bit29 net70 net96 VGND VGND VPWR VPWR ConfigBits\[251\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1042_ W_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0484_ sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1111_ D1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0528_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame4_bit9 net80 net95 VGND VGND VPWR VPWR ConfigBits\[263\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2 net226
+ AD0 AD2 AD3 ConfigBits\[258\] ConfigBits\[259\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0757_ Inst_RegFile_32x4/_0200_ Inst_RegFile_32x4/_0206_ Inst_RegFile_32x4/_0215_
+ Inst_RegFile_32x4/_0221_ A_ADR3 A_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0222_
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0826_ Inst_RegFile_32x4/_0286_ VGND VGND VPWR VPWR AD1 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0688_ Inst_RegFile_32x4__1360_/Q Inst_RegFile_32x4__1396_/Q Inst_RegFile_32x4/_0153_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0154_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1309_ Inst_RegFile_32x4/_0479_ Inst_RegFile_32x4__1462_/Q Inst_RegFile_32x4/_0642_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 JW2BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame1_bit24 net65 net92 VGND VGND VPWR VPWR ConfigBits\[374\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame1_bit13 net53 net92 VGND VGND VPWR VPWR ConfigBits\[363\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1 net21
+ net161 net198 net214 ConfigBits\[298\] ConfigBits\[299\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XW6END_inbuf_3__0_ net233 VGND VGND VPWR VPWR W6BEG_i\[3\] sky130_fd_sc_hd__clkbuf_2
XNN4END_inbuf_7__0_ net139 VGND VGND VPWR VPWR NN4BEG_i\[7\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XEE4BEG_outbuf_0__0_ EE4BEG_i\[0\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1025_ W_ADR4 W_ADR3 W_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0471_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0809_ Inst_RegFile_32x4/_0168_ Inst_RegFile_32x4/_0271_ Inst_RegFile_32x4/_0158_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0272_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput100 FrameStrobe[9] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_16
Xinput133 N4END[6] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput111 N2END[6] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_4
Xinput122 N4END[10] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
Xinput144 NN4END[1] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_4
Xinput199 SS4END[4] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
Xinput177 S4END[13] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xinput188 S4END[9] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
Xinput166 S2MID[1] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_2
Xinput155 S1END[2] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame4_bit28 net69 net95 VGND VGND VPWR VPWR ConfigBits\[282\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame4_bit17 net57 net95 VGND VGND VPWR VPWR ConfigBits\[271\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame11_bit8 net79 net83 VGND VGND VPWR VPWR ConfigBits\[38\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1008_ Inst_RegFile_32x4/_0456_ W_ADR0 Inst_RegFile_32x4/_0457_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0458_ sky130_fd_sc_hd__and3b_2
XFILLER_0_63_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__buf_1
XInst_RegFile_ConfigMem_Inst_frame0_bit12 net52 net81 VGND VGND VPWR VPWR ConfigBits\[394\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame0_bit23 net64 net81 VGND VGND VPWR VPWR ConfigBits\[405\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst1 BD3 J2MID_EFb_BEG\[1\]
+ J2MID_GHb_BEG\[1\] J2END_CD_BEG\[1\] ConfigBits\[24\] ConfigBits\[25\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame0_bit1 net60 net81 VGND VGND VPWR VPWR ConfigBits\[383\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput404 net404 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1 AD0 AD1
+ AD2 AD3 ConfigBits\[50\] ConfigBits\[51\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1290_ Inst_RegFile_32x4/_0634_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0105_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput448 net448 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput437 net437 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput426 net426 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput415 net415 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput459 net459 VGND VGND VPWR VPWR W1BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG1 net115 net167 net220
+ JE2BEG\[6\] ConfigBits\[184\] ConfigBits\[185\] VGND VGND VPWR VPWR J2MID_GHa_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame3_bit16 net56 net94 VGND VGND VPWR VPWR ConfigBits\[302\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix__58_ net220 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1 net153
+ net155 net163 net208 ConfigBits\[370\] ConfigBits\[371\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame3_bit27 net68 net94 VGND VGND VPWR VPWR ConfigBits\[313\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XEE4BEG_outbuf_10__0_ EE4BEG_i\[10\] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0790_ Inst_RegFile_32x4/_0253_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1386_/D
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1342_ net205 Inst_RegFile_32x4/_0002_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1342_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1411_ net205 Inst_RegFile_32x4/_0063_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1411_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput278 net278 VGND VGND VPWR VPWR E6BEG[2] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1273_ Inst_RegFile_32x4/_0624_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0098_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput289 net289 VGND VGND VPWR VPWR EE4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput267 net267 VGND VGND VPWR VPWR E2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput256 net256 VGND VGND VPWR VPWR E1BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG3 net145 net6 net158 net211
+ ConfigBits\[244\] ConfigBits\[245\] VGND VGND VPWR VPWR J2END_EF_BEG\[3\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame7_bit7 net78 net98 VGND VGND VPWR VPWR ConfigBits\[165\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0988_ Inst_RegFile_32x4/_0296_ Inst_RegFile_32x4/_0439_ Inst_RegFile_32x4/_0309_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0440_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0 net101
+ net105 net137 net1 ConfigBits\[282\] ConfigBits\[283\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_23__0_ net64 VGND VGND VPWR VPWR FrameData_O_i\[23\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0911_ Inst_RegFile_32x4__1345_/Q Inst_RegFile_32x4__1393_/Q Inst_RegFile_32x4__1465_/Q
+ Inst_RegFile_32x4__1461_/Q Inst_RegFile_32x4/_0307_ Inst_RegFile_32x4/_0322_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0367_ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0842_ B_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0300_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0773_ Inst_RegFile_32x4/_0233_ Inst_RegFile_32x4/_0235_ Inst_RegFile_32x4/_0236_
+ Inst_RegFile_32x4/_0149_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0237_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_ConfigMem_Inst_frame2_bit26 net67 net93 VGND VGND VPWR VPWR ConfigBits\[344\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst0 net101
+ net1 net206 AD3 ConfigBits\[80\] ConfigBits\[81\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1325_ Inst_RegFile_32x4/_0477_ Inst_RegFile_32x4__1469_/Q Inst_RegFile_32x4/_0652_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0654_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame2_bit15 net55 net93 VGND VGND VPWR VPWR ConfigBits\[333\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1256_ Inst_RegFile_32x4/_0584_ Inst_RegFile_32x4__1439_/Q Inst_RegFile_32x4/_0611_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0615_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1187_ Inst_RegFile_32x4/_0451_ Inst_RegFile_32x4__1412_/Q Inst_RegFile_32x4/_0572_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0573_ sky130_fd_sc_hd__mux2_1
Xstrobe_inbuf_2__0_ net93 VGND VGND VPWR VPWR FrameStrobe_O_i\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_14__0_ net54 VGND VGND VPWR VPWR FrameData_O_i\[14\] sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1 net154
+ net162 net198 net207 ConfigBits\[334\] ConfigBits\[335\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1110_ Inst_RegFile_32x4/_0527_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0032_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XWW4BEG_outbuf_11__0_ WW4BEG_i\[11\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame5_bit19 net59 net96 VGND VGND VPWR VPWR ConfigBits\[241\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1041_ Inst_RegFile_32x4/_0452_ Inst_RegFile_32x4/_0454_ Inst_RegFile_32x4/_0453_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0483_ sky130_fd_sc_hd__or3b_4
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[258\] ConfigBits\[259\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0687_ A_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0153_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0825_ Inst_RegFile_32x4__1385_/D Inst_RegFile_32x4__1385_/Q ConfigBits\[0\]
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0286_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0756_ Inst_RegFile_32x4/_0217_ Inst_RegFile_32x4/_0219_ Inst_RegFile_32x4/_0220_
+ Inst_RegFile_32x4/_0163_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0221_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1239_ Inst_RegFile_32x4/_0605_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0083_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1308_ Inst_RegFile_32x4/_0644_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0113_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 JW2BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_17__0_ FrameStrobe_O_i\[17\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame1_bit25 net66 net92 VGND VGND VPWR VPWR ConfigBits\[375\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame1_bit14 net54 net92 VGND VGND VPWR VPWR ConfigBits\[364\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2 net226
+ AD0 AD1 AD2 ConfigBits\[298\] ConfigBits\[299\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1024_ D0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0470_ sky130_fd_sc_hd__buf_1
XFILLER_0_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0808_ Inst_RegFile_32x4__1451_/Q Inst_RegFile_32x4__1475_/Q Inst_RegFile_32x4/_0156_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0739_ Inst_RegFile_32x4/_0141_ Inst_RegFile_32x4/_0203_ Inst_RegFile_32x4/_0158_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0204_ sky130_fd_sc_hd__a21o_1
Xinput178 S4END[14] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xinput156 S1END[3] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xinput167 S2MID[2] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_2
XWW4END_inbuf_8__0_ net241 VGND VGND VPWR VPWR WW4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_2
Xinput134 N4END[7] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xinput101 N1END[0] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_4
Xinput112 N2END[7] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_4
Xinput123 N4END[11] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput145 NN4END[2] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_2
Xinput189 SS4END[0] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame4_bit29 net70 net95 VGND VGND VPWR VPWR ConfigBits\[283\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame4_bit18 net58 net95 VGND VGND VPWR VPWR ConfigBits\[272\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame11_bit9 net80 net83 VGND VGND VPWR VPWR ConfigBits\[39\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1007_ W_en VGND VGND VPWR VPWR Inst_RegFile_32x4/_0457_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG0 net8 net198 net246 JN2BEG\[2\]
+ ConfigBits\[390\] ConfigBits\[391\] VGND VGND VPWR VPWR J_l_CD_BEG\[0\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame0_bit24 net65 net81 VGND VGND VPWR VPWR ConfigBits\[406\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__1_/A1 ConfigBits\[43\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame0_bit13 net53 net81 VGND VGND VPWR VPWR ConfigBits\[395\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput405 net405 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
XInst_RegFile_ConfigMem_Inst_frame0_bit2 net71 net81 VGND VGND VPWR VPWR ConfigBits\[384\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput416 net416 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2 BD0 BD1
+ BD2 BD3 ConfigBits\[50\] ConfigBits\[51\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput449 net449 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput427 net427 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput438 net438 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG2 net17 net169 net222
+ JS2BEG\[6\] ConfigBits\[186\] ConfigBits\[187\] VGND VGND VPWR VPWR J2MID_GHa_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_70_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame3_bit17 net57 net94 VGND VGND VPWR VPWR ConfigBits\[303\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit28 net69 net94 VGND VGND VPWR VPWR ConfigBits\[314\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__57_ net219 VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2 net246
+ AD0 AD1 AD2 ConfigBits\[370\] ConfigBits\[371\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xstrobe_inbuf_14__0_ net86 VGND VGND VPWR VPWR FrameStrobe_O_i\[14\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XE6END_inbuf_8__0_ net22 VGND VGND VPWR VPWR E6BEG_i\[8\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1272_ Inst_RegFile_32x4__1446_/Q Inst_RegFile_32x4/_0596_ Inst_RegFile_32x4/_0621_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput268 net268 VGND VGND VPWR VPWR E2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput257 net257 VGND VGND VPWR VPWR E1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1410_ net205 Inst_RegFile_32x4/_0062_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1410_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1341_ net205 Inst_RegFile_32x4/_0001_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1341_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput279 net279 VGND VGND VPWR VPWR E6BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame7_bit8 net79 net98 VGND VGND VPWR VPWR ConfigBits\[166\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0987_ Inst_RegFile_32x4__1435_/Q Inst_RegFile_32x4__1431_/Q Inst_RegFile_32x4/_0298_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1 net5 net153
+ net157 net206 ConfigBits\[282\] ConfigBits\[283\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XE6BEG_outbuf_0__0_ E6BEG_i\[0\] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0841_ Inst_RegFile_32x4__1404_/Q Inst_RegFile_32x4__1380_/Q Inst_RegFile_32x4/_0298_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0299_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0910_ Inst_RegFile_32x4/_0302_ Inst_RegFile_32x4/_0365_ Inst_RegFile_32x4/_0319_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0366_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame2_bit27 net68 net93 VGND VGND VPWR VPWR ConfigBits\[345\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame2_bit16 net56 net93 VGND VGND VPWR VPWR ConfigBits\[334\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0772_ Inst_RegFile_32x4__1346_/Q Inst_RegFile_32x4__1394_/Q Inst_RegFile_32x4__1466_/Q
+ Inst_RegFile_32x4__1462_/Q Inst_RegFile_32x4/_0146_ Inst_RegFile_32x4/_0161_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0236_ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1255_ Inst_RegFile_32x4/_0614_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0090_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst1 BD3 J2MID_EFb_BEG\[1\]
+ J2MID_GHb_BEG\[1\] J2END_CD_BEG\[3\] ConfigBits\[80\] ConfigBits\[81\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1324_ Inst_RegFile_32x4/_0653_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0120_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1186_ Inst_RegFile_32x4/_0570_ Inst_RegFile_32x4/_0571_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0572_ sky130_fd_sc_hd__nand2_2
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2 net209
+ AD0 AD1 AD2 ConfigBits\[334\] ConfigBits\[335\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XEE4END_inbuf_9__0_ net37 VGND VGND VPWR VPWR EE4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_2
Xdata_inbuf_6__0_ net77 VGND VGND VPWR VPWR FrameData_O_i\[6\] sky130_fd_sc_hd__buf_1
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1040_ Inst_RegFile_32x4/_0482_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0007_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__1_/A1 ConfigBits\[26\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0824_ Inst_RegFile_32x4/_0285_ VGND VGND VPWR VPWR AD0 sky130_fd_sc_hd__buf_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3/X ConfigBits\[260\]
+ ConfigBits\[261\] VGND VGND VPWR VPWR JN2BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0686_ Inst_RegFile_32x4/_0128_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0152_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0755_ Inst_RegFile_32x4__1409_/Q Inst_RegFile_32x4__1341_/Q Inst_RegFile_32x4__1401_/Q
+ Inst_RegFile_32x4__1469_/Q Inst_RegFile_32x4/_0160_ Inst_RegFile_32x4/_0188_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0220_ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1238_ Inst_RegFile_32x4/_0584_ Inst_RegFile_32x4__1431_/Q Inst_RegFile_32x4/_0601_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0605_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1307_ Inst_RegFile_32x4/_0477_ Inst_RegFile_32x4__1461_/Q Inst_RegFile_32x4/_0642_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0644_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1169_ Inst_RegFile_32x4__1405_/Q Inst_RegFile_32x4/_0528_ Inst_RegFile_32x4/_0560_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 JW2BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame1_bit15 net55 net92 VGND VGND VPWR VPWR ConfigBits\[365\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame1_bit26 net67 net92 VGND VGND VPWR VPWR ConfigBits\[376\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit0 net49 net94 VGND VGND VPWR VPWR ConfigBits\[286\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[298\] ConfigBits\[299\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1023_ Inst_RegFile_32x4/_0469_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0003_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0807_ Inst_RegFile_32x4/_0152_ Inst_RegFile_32x4/_0269_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0270_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0738_ Inst_RegFile_32x4__1353_/Q Inst_RegFile_32x4__1349_/Q Inst_RegFile_32x4/_0156_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0669_ Inst_RegFile_32x4/_0134_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0135_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput179 S4END[15] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
Xinput168 S2MID[3] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
Xinput157 S2END[0] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_4
Xinput102 N1END[1] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_4
Xinput113 N2MID[0] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
Xinput135 N4END[8] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
Xinput124 N4END[12] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
Xinput146 NN4END[3] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame4_bit19 net59 net95 VGND VGND VPWR VPWR ConfigBits\[273\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XNN4BEG_outbuf_0__0_ NN4BEG_i\[0\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4BEG_outbuf_4__0_ N4BEG_i\[4\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1006_ W_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0456_ sky130_fd_sc_hd__clkbuf_2
XSS4BEG_outbuf_3__0_ SS4BEG_i\[3\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG1 net129 net7 net217 JE2BEG\[2\]
+ ConfigBits\[392\] ConfigBits\[393\] VGND VGND VPWR VPWR J_l_CD_BEG\[1\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame0_bit25 net66 net81 VGND VGND VPWR VPWR ConfigBits\[407\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame0_bit14 net54 net81 VGND VGND VPWR VPWR ConfigBits\[396\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XSS4BEG_outbuf_11__0_ SS4BEG_i\[11\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame0_bit3 net74 net81 VGND VGND VPWR VPWR ConfigBits\[385\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3 J2MID_ABb_BEG\[1\]
+ J2MID_CDb_BEG\[1\] J2MID_EFb_BEG\[1\] J2MID_GHb_BEG\[1\] ConfigBits\[50\] ConfigBits\[51\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput428 net428 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput439 net439 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput417 net417 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput406 net406 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XW6BEG_outbuf_4__0_ W6BEG_i\[4\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG3 net113 net13 net218
+ JW2BEG\[6\] ConfigBits\[188\] ConfigBits\[189\] VGND VGND VPWR VPWR J2MID_GHa_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame3_bit18 net58 net94 VGND VGND VPWR VPWR ConfigBits\[304\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit29 net70 net94 VGND VGND VPWR VPWR ConfigBits\[315\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__56_ net218 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3 AD3 BD0
+ BD2 BD3 ConfigBits\[370\] ConfigBits\[371\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__1_/A1 ConfigBits\[105\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1271_ Inst_RegFile_32x4/_0623_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0097_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput269 net269 VGND VGND VPWR VPWR E2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput258 net258 VGND VGND VPWR VPWR E2BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1340_ net205 Inst_RegFile_32x4/_0000_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1340_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame7_bit9 net80 net98 VGND VGND VPWR VPWR ConfigBits\[167\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0986_ Inst_RegFile_32x4/_0290_ Inst_RegFile_32x4/_0437_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0438_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_24__0_ FrameData_O_i\[24\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2 net208
+ AD0 AD1 AD2 ConfigBits\[282\] ConfigBits\[283\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1469_ net205 Inst_RegFile_32x4/_0121_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1469_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__39_ JS2BEG\[7\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_outbuf_15__0_ FrameData_O_i\[15\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_4__0_ S4BEG_i\[4\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0840_ Inst_RegFile_32x4/_0297_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0298_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0771_ Inst_RegFile_32x4/_0141_ Inst_RegFile_32x4/_0234_ Inst_RegFile_32x4/_0158_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame2_bit17 net57 net93 VGND VGND VPWR VPWR ConfigBits\[335\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame2_bit28 net69 net93 VGND VGND VPWR VPWR ConfigBits\[346\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1254_ Inst_RegFile_32x4/_0582_ Inst_RegFile_32x4__1438_/Q Inst_RegFile_32x4/_0611_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0614_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1185_ W_ADR2 W_ADR3 W_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0571_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1323_ Inst_RegFile_32x4/_0470_ Inst_RegFile_32x4__1468_/Q Inst_RegFile_32x4/_0652_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3 AD3 BD1
+ BD2 BD3 ConfigBits\[334\] ConfigBits\[335\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0969_ Inst_RegFile_32x4/_0346_ Inst_RegFile_32x4/_0420_ Inst_RegFile_32x4/_0300_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XS4END_inbuf_2__0_ net185 VGND VGND VPWR VPWR S4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0754_ Inst_RegFile_32x4/_0185_ Inst_RegFile_32x4/_0218_ Inst_RegFile_32x4/_0171_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0219_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0823_ Inst_RegFile_32x4__1384_/D Inst_RegFile_32x4__1384_/Q ConfigBits\[0\]
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XEE4BEG_outbuf_3__0_ EE4BEG_i\[3\] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0685_ Inst_RegFile_32x4/_0133_ Inst_RegFile_32x4/_0140_ Inst_RegFile_32x4/_0144_
+ Inst_RegFile_32x4/_0150_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0151_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XW6END_inbuf_6__0_ net236 VGND VGND VPWR VPWR W6BEG_i\[6\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1306_ Inst_RegFile_32x4/_0643_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0112_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1237_ Inst_RegFile_32x4/_0604_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0082_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1168_ Inst_RegFile_32x4/_0561_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0056_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1099_ Inst_RegFile_32x4/_0520_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0028_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame1_bit27 net68 net92 VGND VGND VPWR VPWR ConfigBits\[377\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame1_bit16 net56 net92 VGND VGND VPWR VPWR ConfigBits\[366\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame3_bit1 net60 net94 VGND VGND VPWR VPWR ConfigBits\[287\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3/X ConfigBits\[300\]
+ ConfigBits\[301\] VGND VGND VPWR VPWR JE2BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1022_ Inst_RegFile_32x4/_0468_ Inst_RegFile_32x4__1343_/Q Inst_RegFile_32x4/_0459_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0469_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0806_ Inst_RegFile_32x4__1459_/Q Inst_RegFile_32x4__1455_/Q Inst_RegFile_32x4/_0153_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0737_ Inst_RegFile_32x4/_0188_ Inst_RegFile_32x4/_0201_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0202_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0668_ A_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0134_ sky130_fd_sc_hd__buf_2
Xinput169 S2MID[4] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_2
Xinput158 S2END[1] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_4
Xinput103 N1END[2] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_4
Xinput114 N2MID[1] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xinput136 N4END[9] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
Xinput125 N4END[13] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
Xinput147 NN4END[4] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0 net104
+ net106 net6 net24 ConfigBits\[350\] ConfigBits\[351\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1005_ Inst_RegFile_32x4/_0452_ Inst_RegFile_32x4/_0453_ Inst_RegFile_32x4/_0454_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0455_ sky130_fd_sc_hd__and3_2
XFILLER_0_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG2 net144 net40 net180 JS2BEG\[2\]
+ ConfigBits\[394\] ConfigBits\[395\] VGND VGND VPWR VPWR J_l_CD_BEG\[2\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame0_bit26 net67 net81 VGND VGND VPWR VPWR ConfigBits\[408\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame0_bit15 net55 net81 VGND VGND VPWR VPWR ConfigBits\[397\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame0_bit4 net75 net81 VGND VGND VPWR VPWR ConfigBits\[386\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3/X ConfigBits\[52\]
+ ConfigBits\[53\] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__mux4_2
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput429 net429 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput418 net418 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput407 net407 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame10_bit0 net49 net82 VGND VGND VPWR VPWR ConfigBits\[62\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XN4END_inbuf_10__0_ net126 VGND VGND VPWR VPWR N4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix__55_ JW2BEG\[7\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame3_bit19 net59 net94 VGND VGND VPWR VPWR ConfigBits\[305\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3/X ConfigBits\[372\]
+ ConfigBits\[373\] VGND VGND VPWR VPWR JW2BEG\[5\] sky130_fd_sc_hd__mux4_2
XFILLER_0_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_2__0_ FrameData_O_i\[2\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1270_ Inst_RegFile_32x4__1445_/Q Inst_RegFile_32x4/_0594_ Inst_RegFile_32x4/_0621_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0623_ sky130_fd_sc_hd__mux2_1
Xoutput259 net259 VGND VGND VPWR VPWR E2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xdata_inbuf_26__0_ net67 VGND VGND VPWR VPWR FrameData_O_i\[26\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0985_ Inst_RegFile_32x4__1443_/Q Inst_RegFile_32x4__1439_/Q Inst_RegFile_32x4/_0335_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0437_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3 AD3 BD0
+ BD1 BD2 ConfigBits\[282\] ConfigBits\[283\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1468_ net205 Inst_RegFile_32x4/_0120_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1468_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xstrobe_inbuf_5__0_ net96 VGND VGND VPWR VPWR FrameStrobe_O_i\[5\] sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix__38_ JS2BEG\[6\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1399_ net205 Inst_RegFile_32x4/_0051_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1399_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xdata_inbuf_17__0_ net57 VGND VGND VPWR VPWR FrameData_O_i\[17\] sky130_fd_sc_hd__buf_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__1_/A1 ConfigBits\[79\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG0 net120 net20 net172
+ net225 ConfigBits\[198\] ConfigBits\[199\] VGND VGND VPWR VPWR J2MID_CDb_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR A_ADR4 sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_E1BEG0 AD3 J2MID_CDb_BEG\[3\] JN2BEG\[3\]
+ J_l_CD_BEG\[1\] ConfigBits\[30\] ConfigBits\[31\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__0770_ Inst_RegFile_32x4__1354_/Q Inst_RegFile_32x4__1350_/Q Inst_RegFile_32x4/_0142_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame2_bit18 net58 net93 VGND VGND VPWR VPWR ConfigBits\[336\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame2_bit29 net70 net93 VGND VGND VPWR VPWR ConfigBits\[347\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1322_ Inst_RegFile_32x4/_0455_ Inst_RegFile_32x4/_0570_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0652_ sky130_fd_sc_hd__nand2_2
XInst_RegFile_32x4__1253_ Inst_RegFile_32x4/_0613_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0089_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1184_ Inst_RegFile_32x4/_0456_ Inst_RegFile_32x4/_0484_ Inst_RegFile_32x4/_0457_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0570_ sky130_fd_sc_hd__and3_2
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3/X ConfigBits\[336\]
+ ConfigBits\[337\] VGND VGND VPWR VPWR JS2BEG\[4\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__0968_ Inst_RegFile_32x4__1407_/Q Inst_RegFile_32x4__1383_/Q Inst_RegFile_32x4/_0298_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0420_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0899_ Inst_RegFile_32x4/_0290_ Inst_RegFile_32x4/_0354_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0355_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4END_inbuf_10__0_ net178 VGND VGND VPWR VPWR S4BEG_i\[10\] sky130_fd_sc_hd__buf_2
XFILLER_0_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0822_ Inst_RegFile_32x4/_0284_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1387_/D
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0753_ Inst_RegFile_32x4__1417_/Q Inst_RegFile_32x4__1413_/Q Inst_RegFile_32x4/_0169_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0218_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0684_ Inst_RegFile_32x4/_0145_ Inst_RegFile_32x4/_0147_ Inst_RegFile_32x4/_0149_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0150_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1305_ Inst_RegFile_32x4/_0470_ Inst_RegFile_32x4__1460_/Q Inst_RegFile_32x4/_0642_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0643_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1236_ Inst_RegFile_32x4/_0582_ Inst_RegFile_32x4__1430_/Q Inst_RegFile_32x4/_0601_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0604_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1167_ Inst_RegFile_32x4__1404_/Q Inst_RegFile_32x4/_0524_ Inst_RegFile_32x4/_0560_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0561_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1098_ Inst_RegFile_32x4__1368_/Q Inst_RegFile_32x4/_0491_ Inst_RegFile_32x4/_0519_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame1_bit17 net57 net92 VGND VGND VPWR VPWR ConfigBits\[367\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame1_bit28 net69 net92 VGND VGND VPWR VPWR ConfigBits\[378\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame3_bit2 net71 net94 VGND VGND VPWR VPWR ConfigBits\[288\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1021_ Inst_RegFile_32x4/_0467_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0468_
+ sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__0667_ Inst_RegFile_32x4/_0129_ Inst_RegFile_32x4/_0132_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0133_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0805_ Inst_RegFile_32x4/_0264_ Inst_RegFile_32x4/_0266_ Inst_RegFile_32x4/_0267_
+ Inst_RegFile_32x4/_0149_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0268_ sky130_fd_sc_hd__o22a_2
XInst_RegFile_32x4__0736_ Inst_RegFile_32x4__1361_/Q Inst_RegFile_32x4__1397_/Q Inst_RegFile_32x4/_0153_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0201_ sky130_fd_sc_hd__mux2_1
XSS4END_inbuf_0__0_ net199 VGND VGND VPWR VPWR SS4BEG_i\[0\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1219_ Inst_RegFile_32x4__1424_/Q Inst_RegFile_32x4/_0591_ Inst_RegFile_32x4/_0592_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0593_ sky130_fd_sc_hd__mux2_1
Xinput115 N2MID[2] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
Xinput104 N1END[3] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_8
Xinput126 N4END[14] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
Xinput159 S2END[2] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
Xinput148 NN4END[5] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xinput137 NN4END[0] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_2__0_ FrameStrobe_O_i\[2\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1 net158
+ net180 net189 net211 ConfigBits\[350\] ConfigBits\[351\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1004_ W_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0454_ sky130_fd_sc_hd__buf_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG3 net121 net189 net226 JW2BEG\[2\]
+ ConfigBits\[396\] ConfigBits\[397\] VGND VGND VPWR VPWR J_l_CD_BEG\[3\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame0_bit16 net56 net81 VGND VGND VPWR VPWR ConfigBits\[398\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0719_ Inst_RegFile_32x4/_0134_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0185_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame0_bit27 net68 net81 VGND VGND VPWR VPWR ConfigBits\[409\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_17__0_ net89 VGND VGND VPWR VPWR FrameStrobe_O_i\[17\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame0_bit5 net76 net81 VGND VGND VPWR VPWR ConfigBits\[387\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XWW4BEG_outbuf_0__0_ WW4BEG_i\[0\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0 net108
+ net130 net2 net8 ConfigBits\[262\] ConfigBits\[263\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
Xoutput419 net419 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput408 net408 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_0_10_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame10_bit1 net60 net82 VGND VGND VPWR VPWR ConfigBits\[63\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_A_ADR0 J2MID_EFa_BEG\[0\] J2MID_EFb_BEG\[0\]
+ J2END_EF_BEG\[0\] J_l_EF_BEG\[0\] ConfigBits\[114\] ConfigBits\[115\] VGND VGND
+ VPWR VPWR A_ADR0 sky130_fd_sc_hd__mux4_2
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix__54_ JW2BEG\[6\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XE6BEG_outbuf_3__0_ E6BEG_i\[3\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG0 net119 net171 net224
+ JN2BEG\[3\] ConfigBits\[158\] ConfigBits\[159\] VGND VGND VPWR VPWR J2MID_ABa_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XN4END_inbuf_2__0_ net133 VGND VGND VPWR VPWR N4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0984_ Inst_RegFile_32x4/_0329_ Inst_RegFile_32x4/_0435_ Inst_RegFile_32x4/_0319_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0436_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3/X ConfigBits\[284\]
+ ConfigBits\[285\] VGND VGND VPWR VPWR JN2BEG\[7\] sky130_fd_sc_hd__mux4_2
XFILLER_0_60_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1467_ net205 Inst_RegFile_32x4/_0119_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1467_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1398_ net205 Inst_RegFile_32x4/_0050_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1398_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__37_ JS2BEG\[5\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame6_bit0 net49 net97 VGND VGND VPWR VPWR ConfigBits\[190\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_9__0_ net80 VGND VGND VPWR VPWR FrameData_O_i\[9\] sky130_fd_sc_hd__buf_1
XFILLER_0_51_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_E1BEG1 BD0 J2MID_EFb_BEG\[0\] JN2BEG\[0\]
+ J_l_EF_BEG\[2\] ConfigBits\[32\] ConfigBits\[33\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__mux4_2
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_my_mux2_inst__1_/A1 ConfigBits\[124\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG1 net116 net16 net168
+ net221 ConfigBits\[200\] ConfigBits\[201\] VGND VGND VPWR VPWR J2MID_CDb_BEG\[1\]
+ sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__1252_ Inst_RegFile_32x4/_0580_ Inst_RegFile_32x4__1437_/Q Inst_RegFile_32x4/_0611_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0613_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame2_bit19 net59 net93 VGND VGND VPWR VPWR ConfigBits\[337\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1321_ Inst_RegFile_32x4/_0651_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0119_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst0 net104
+ net4 net156 AD2 ConfigBits\[41\] ConfigBits\[42\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1183_ Inst_RegFile_32x4/_0569_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0063_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0967_ Inst_RegFile_32x4/_0343_ Inst_RegFile_32x4/_0418_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0419_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0898_ Inst_RegFile_32x4__1357_/Q Inst_RegFile_32x4__1445_/Q Inst_RegFile_32x4/_0292_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0821_ Inst_RegFile_32x4/_0262_ Inst_RegFile_32x4/_0268_ Inst_RegFile_32x4/_0277_
+ Inst_RegFile_32x4/_0283_ A_ADR3 A_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0284_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0752_ Inst_RegFile_32x4/_0182_ Inst_RegFile_32x4/_0216_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0217_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0683_ Inst_RegFile_32x4/_0148_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0149_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1235_ Inst_RegFile_32x4/_0603_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0081_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1304_ Inst_RegFile_32x4/_0471_ Inst_RegFile_32x4/_0570_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0642_ sky130_fd_sc_hd__nand2_2
XInst_RegFile_32x4__1166_ Inst_RegFile_32x4/_0493_ Inst_RegFile_32x4/_0502_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0560_ sky130_fd_sc_hd__nor2_2
XInst_RegFile_32x4__1097_ Inst_RegFile_32x4/_0493_ Inst_RegFile_32x4/_0513_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0519_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame1_bit29 net70 net92 VGND VGND VPWR VPWR ConfigBits\[379\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame1_bit18 net58 net92 VGND VGND VPWR VPWR ConfigBits\[368\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame3_bit3 net74 net94 VGND VGND VPWR VPWR ConfigBits\[289\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XNN4BEG_outbuf_3__0_ NN4BEG_i\[3\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1020_ D3 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0467_ sky130_fd_sc_hd__clkbuf_2
XN4BEG_outbuf_7__0_ N4BEG_i\[7\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0804_ Inst_RegFile_32x4__1347_/Q Inst_RegFile_32x4__1395_/Q Inst_RegFile_32x4__1467_/Q
+ Inst_RegFile_32x4__1463_/Q Inst_RegFile_32x4/_0146_ Inst_RegFile_32x4/_0134_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0267_ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0666_ Inst_RegFile_32x4__1356_/Q Inst_RegFile_32x4__1444_/Q Inst_RegFile_32x4/_0131_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0735_ Inst_RegFile_32x4/_0193_ Inst_RegFile_32x4/_0195_ Inst_RegFile_32x4/_0197_
+ Inst_RegFile_32x4/_0199_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0200_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_32x4__1218_ Inst_RegFile_32x4/_0474_ Inst_RegFile_32x4/_0571_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0592_ sky130_fd_sc_hd__and2_2
Xinput138 NN4END[10] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
XSS4BEG_outbuf_6__0_ SS4BEG_i\[6\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_1
Xinput116 N2MID[3] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput105 N2END[0] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_4
Xinput149 NN4END[6] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
Xinput127 N4END[15] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1149_ Inst_RegFile_32x4/_0550_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0048_
+ sky130_fd_sc_hd__clkbuf_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XS4BEG_outbuf_10__0_ S4BEG_i\[10\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2 net229
+ AD1 AD2 AD3 ConfigBits\[350\] ConfigBits\[351\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XW6BEG_outbuf_7__0_ W6BEG_i\[7\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1003_ W_ADR3 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0453_ sky130_fd_sc_hd__buf_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0718_ Inst_RegFile_32x4/_0182_ Inst_RegFile_32x4/_0183_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0184_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame0_bit17 net57 net81 VGND VGND VPWR VPWR ConfigBits\[399\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame0_bit28 net69 net81 VGND VGND VPWR VPWR ConfigBits\[410\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame0_bit6 net77 net81 VGND VGND VPWR VPWR ConfigBits\[388\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1 net24
+ net160 net213 net246 ConfigBits\[262\] ConfigBits\[263\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xoutput409 net409 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XNN4END_inbuf_0__0_ net147 VGND VGND VPWR VPWR NN4BEG_i\[0\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame10_bit2 net71 net82 VGND VGND VPWR VPWR ConfigBits\[64\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_A_ADR1 J2MID_EFa_BEG\[1\] J2MID_EFb_BEG\[1\]
+ J2END_EF_BEG\[1\] J_l_EF_BEG\[1\] ConfigBits\[116\] ConfigBits\[117\] VGND VGND
+ VPWR VPWR A_ADR1 sky130_fd_sc_hd__mux4_2
XFILLER_0_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__53_ JW2BEG\[5\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_27__0_ FrameData_O_i\[27\] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0 net102
+ net110 net2 net10 ConfigBits\[302\] ConfigBits\[303\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_outbuf_18__0_ FrameData_O_i\[18\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG1 net15 net167 net220
+ JE2BEG\[3\] ConfigBits\[160\] ConfigBits\[161\] VGND VGND VPWR VPWR J2MID_ABa_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XS4BEG_outbuf_7__0_ S4BEG_i\[7\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0983_ Inst_RegFile_32x4__1451_/Q Inst_RegFile_32x4__1475_/Q Inst_RegFile_32x4/_0317_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1397_ net205 Inst_RegFile_32x4/_0049_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1397_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1466_ net205 Inst_RegFile_32x4/_0118_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1466_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__36_ JS2BEG\[4\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XS4END_inbuf_5__0_ net188 VGND VGND VPWR VPWR S4BEG_i\[5\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame6_bit1 net60 net97 VGND VGND VPWR VPWR ConfigBits\[191\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_E1BEG2 BD1 J2MID_GHb_BEG\[1\] JN2BEG\[1\]
+ J_l_GH_BEG\[3\] ConfigBits\[34\] ConfigBits\[35\] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG2 net118 net18 net170
+ net223 ConfigBits\[202\] ConfigBits\[203\] VGND VGND VPWR VPWR J2MID_CDb_BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1251_ Inst_RegFile_32x4/_0612_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0088_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1182_ Inst_RegFile_32x4/_0468_ Inst_RegFile_32x4__1411_/Q Inst_RegFile_32x4/_0565_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0569_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1320_ Inst_RegFile_32x4/_0481_ Inst_RegFile_32x4__1467_/Q Inst_RegFile_32x4/_0647_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0651_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst1 BD2 J2MID_ABa_BEG\[2\]
+ J2MID_CDa_BEG\[2\] J2END_EF_BEG\[0\] ConfigBits\[41\] ConfigBits\[42\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0966_ Inst_RegFile_32x4__1359_/Q Inst_RegFile_32x4__1447_/Q Inst_RegFile_32x4/_0292_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0418_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0897_ Inst_RegFile_32x4/_0353_ VGND VGND VPWR VPWR BD0 sky130_fd_sc_hd__buf_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst0 net102
+ net2 net207 AD0 ConfigBits\[27\] ConfigBits\[28\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XEE4BEG_outbuf_6__0_ EE4BEG_i\[6\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XW6END_inbuf_9__0_ net228 VGND VGND VPWR VPWR W6BEG_i\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1449_ net205 Inst_RegFile_32x4/_0101_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1449_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__19_ JN2BEG\[3\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0 net146
+ net3 net198 net208 ConfigBits\[54\] ConfigBits\[55\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0751_ Inst_RegFile_32x4__1425_/Q Inst_RegFile_32x4__1421_/Q Inst_RegFile_32x4/_0165_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0216_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0820_ Inst_RegFile_32x4/_0279_ Inst_RegFile_32x4/_0281_ Inst_RegFile_32x4/_0282_
+ Inst_RegFile_32x4/_0163_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0283_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0682_ A_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0148_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1303_ Inst_RegFile_32x4/_0641_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0111_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1234_ Inst_RegFile_32x4/_0580_ Inst_RegFile_32x4__1429_/Q Inst_RegFile_32x4/_0601_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0603_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0 net104
+ net112 net4 net12 ConfigBits\[374\] ConfigBits\[375\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1165_ Inst_RegFile_32x4/_0559_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0055_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1096_ Inst_RegFile_32x4/_0518_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0027_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0949_ Inst_RegFile_32x4__1450_/Q Inst_RegFile_32x4__1474_/Q Inst_RegFile_32x4/_0317_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame1_bit19 net59 net92 VGND VGND VPWR VPWR ConfigBits\[369\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame3_bit4 net75 net94 VGND VGND VPWR VPWR ConfigBits\[290\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0734_ Inst_RegFile_32x4/_0145_ Inst_RegFile_32x4/_0198_ Inst_RegFile_32x4/_0149_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0199_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0803_ Inst_RegFile_32x4/_0141_ Inst_RegFile_32x4/_0265_ A_ADR2
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0266_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0665_ Inst_RegFile_32x4/_0130_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0131_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1217_ D0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0591_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1148_ Inst_RegFile_32x4__1396_/Q Inst_RegFile_32x4/_0524_ Inst_RegFile_32x4/_0549_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0550_ sky130_fd_sc_hd__mux2_1
Xinput139 NN4END[11] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xinput117 N2MID[4] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
Xinput106 N2END[1] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
Xinput128 N4END[1] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1079_ Inst_RegFile_32x4__1360_/Q Inst_RegFile_32x4/_0491_ Inst_RegFile_32x4/_0508_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0509_ sky130_fd_sc_hd__mux2_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XNN4BEG_outbuf_10__0_ NN4BEG_i\[10\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[350\] ConfigBits\[351\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0 net103
+ net111 net3 net11 ConfigBits\[338\] ConfigBits\[339\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1002_ W_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0452_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0717_ Inst_RegFile_32x4__1424_/Q Inst_RegFile_32x4__1420_/Q Inst_RegFile_32x4/_0131_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame0_bit18 net58 net81 VGND VGND VPWR VPWR ConfigBits\[400\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame0_bit29 net70 net81 VGND VGND VPWR VPWR ConfigBits\[411\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame0_bit7 net78 net81 VGND VGND VPWR VPWR ConfigBits\[389\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_outbuf_10__0_ FrameStrobe_O_i\[10\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_outbuf_5__0_ FrameData_O_i\[5\] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2 net229
+ AD0 AD1 AD3 ConfigBits\[262\] ConfigBits\[263\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame10_bit3 net74 net82 VGND VGND VPWR VPWR ConfigBits\[65\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_A_ADR2 J2MID_EFa_BEG\[2\] J2MID_EFb_BEG\[2\]
+ J2END_EF_BEG\[2\] J_l_EF_BEG\[2\] ConfigBits\[118\] ConfigBits\[119\] VGND VGND
+ VPWR VPWR A_ADR2 sky130_fd_sc_hd__mux4_2
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_29__0_ net70 VGND VGND VPWR VPWR FrameData_O_i\[29\] sky130_fd_sc_hd__clkbuf_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__52_ JW2BEG\[4\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XWW4END_inbuf_1__0_ net249 VGND VGND VPWR VPWR WW4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_8__0_ net99 VGND VGND VPWR VPWR FrameStrobe_O_i\[8\] sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1 net42
+ net154 net156 net162 ConfigBits\[302\] ConfigBits\[303\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG2 net117 net17 net222
+ JS2BEG\[3\] ConfigBits\[162\] ConfigBits\[163\] VGND VGND VPWR VPWR J2MID_ABa_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0982_ Inst_RegFile_32x4/_0313_ Inst_RegFile_32x4/_0433_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0434_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1396_ net205 Inst_RegFile_32x4/_0048_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1396_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__35_ JS2BEG\[3\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1465_ net205 Inst_RegFile_32x4/_0117_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1465_/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame6_bit2 net71 net97 VGND VGND VPWR VPWR ConfigBits\[192\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_E1BEG3 BD2 J2MID_ABb_BEG\[2\] JN2BEG\[2\]
+ J_l_AB_BEG\[0\] ConfigBits\[36\] ConfigBits\[37\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__mux4_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG3 net114 net14 net166
+ net219 ConfigBits\[204\] ConfigBits\[205\] VGND VGND VPWR VPWR J2MID_CDb_BEG\[3\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1250_ Inst_RegFile_32x4/_0577_ Inst_RegFile_32x4__1436_/Q Inst_RegFile_32x4/_0611_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1181_ Inst_RegFile_32x4/_0568_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0062_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0965_ Inst_RegFile_32x4/_0417_ VGND VGND VPWR VPWR BD2 sky130_fd_sc_hd__buf_12
XInst_RegFile_32x4__0896_ Inst_RegFile_32x4__1388_/D Inst_RegFile_32x4__1388_/Q ConfigBits\[1\]
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0353_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR W_en sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1448_ net205 Inst_RegFile_32x4/_0100_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1448_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst1 BD0 J2MID_EFa_BEG\[2\]
+ J2MID_GHa_BEG\[2\] J2END_AB_BEG\[1\] ConfigBits\[27\] ConfigBits\[28\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix__18_ JN2BEG\[2\] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__1379_ net205 Inst_RegFile_32x4/_0039_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1379_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1 AD0 AD1
+ AD2 AD3 ConfigBits\[54\] ConfigBits\[55\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XE6END_inbuf_1__0_ net26 VGND VGND VPWR VPWR E6BEG_i\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0750_ Inst_RegFile_32x4/_0208_ Inst_RegFile_32x4/_0210_ Inst_RegFile_32x4/_0212_
+ Inst_RegFile_32x4/_0214_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0215_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1302_ Inst_RegFile_32x4__1459_/Q Inst_RegFile_32x4/_0467_ Inst_RegFile_32x4/_0637_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0641_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0681_ Inst_RegFile_32x4__1368_/Q Inst_RegFile_32x4__1364_/Q Inst_RegFile_32x4/_0146_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1 net154
+ net156 net164 net209 ConfigBits\[374\] ConfigBits\[375\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1233_ Inst_RegFile_32x4/_0602_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0080_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1095_ Inst_RegFile_32x4__1367_/Q Inst_RegFile_32x4/_0500_ Inst_RegFile_32x4/_0514_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0518_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1164_ Inst_RegFile_32x4/_0468_ Inst_RegFile_32x4__1403_/Q Inst_RegFile_32x4/_0555_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0559_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0948_ Inst_RegFile_32x4/_0313_ Inst_RegFile_32x4/_0401_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0402_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0879_ Inst_RegFile_32x4/_0334_ Inst_RegFile_32x4/_0336_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0337_ sky130_fd_sc_hd__and2b_1
XSS4END_inbuf_3__0_ net202 VGND VGND VPWR VPWR SS4BEG_i\[3\] sky130_fd_sc_hd__buf_2
XFILLER_0_61_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput390 net390 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame3_bit5 net76 net94 VGND VGND VPWR VPWR ConfigBits\[291\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_5__0_ FrameStrobe_O_i\[5\] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0664_ A_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0130_ sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__0733_ Inst_RegFile_32x4__1369_/Q Inst_RegFile_32x4__1365_/Q Inst_RegFile_32x4/_0146_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0802_ Inst_RegFile_32x4__1355_/Q Inst_RegFile_32x4__1351_/Q Inst_RegFile_32x4/_0142_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1216_ Inst_RegFile_32x4/_0590_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0075_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1147_ Inst_RegFile_32x4/_0525_ Inst_RegFile_32x4/_0483_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0549_ sky130_fd_sc_hd__nor2_2
XInst_RegFile_32x4__1078_ Inst_RegFile_32x4/_0473_ Inst_RegFile_32x4/_0483_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0508_ sky130_fd_sc_hd__nor2_2
Xinput118 N2MID[5] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_2
Xinput107 N2END[2] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_4
Xinput129 N4END[2] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XEE4END_inbuf_2__0_ net45 VGND VGND VPWR VPWR EE4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst0 net102
+ net2 net207 AD0 ConfigBits\[83\] ConfigBits\[84\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3/X ConfigBits\[352\]
+ ConfigBits\[353\] VGND VGND VPWR VPWR JW2BEG\[0\] sky130_fd_sc_hd__mux4_2
XFILLER_0_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XWW4BEG_outbuf_3__0_ WW4BEG_i\[3\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__clkbuf_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1 net155
+ net163 net197 net206 ConfigBits\[338\] ConfigBits\[339\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1001_ Inst_RegFile_32x4/_0450_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0451_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0716_ Inst_RegFile_32x4/_0128_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0182_
+ sky130_fd_sc_hd__buf_1
XFILLER_0_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame0_bit19 net59 net81 VGND VGND VPWR VPWR ConfigBits\[401\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame0_bit8 net79 net81 VGND VGND VPWR VPWR ConfigBits\[390\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XE6BEG_outbuf_6__0_ E6BEG_i\[6\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[262\] ConfigBits\[263\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame9_bit0 net49 net100 VGND VGND VPWR VPWR ConfigBits\[94\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit4 net75 net82 VGND VGND VPWR VPWR ConfigBits\[66\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XN4END_inbuf_5__0_ net136 VGND VGND VPWR VPWR N4BEG_i\[5\] sky130_fd_sc_hd__buf_2
XInst_RegFile_switch_matrix__51_ JW2BEG\[3\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_A_ADR3 J2MID_EFa_BEG\[3\] J2MID_EFb_BEG\[3\]
+ J2END_EF_BEG\[3\] J_l_EF_BEG\[3\] ConfigBits\[120\] ConfigBits\[121\] VGND VGND
+ VPWR VPWR A_ADR3 sky130_fd_sc_hd__mux4_2
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2 net207
+ AD0 AD1 AD2 ConfigBits\[302\] ConfigBits\[303\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG3 net113 net13 net165
+ JW2BEG\[3\] ConfigBits\[164\] ConfigBits\[165\] VGND VGND VPWR VPWR J2MID_ABa_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0981_ Inst_RegFile_32x4__1459_/Q Inst_RegFile_32x4__1455_/Q Inst_RegFile_32x4/_0314_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1464_ net205 Inst_RegFile_32x4/_0116_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1464_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__34_ JS2BEG\[2\] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1395_ net205 Inst_RegFile_32x4/_0047_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1395_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame6_bit3 net74 net97 VGND VGND VPWR VPWR ConfigBits\[193\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1180_ Inst_RegFile_32x4/_0465_ Inst_RegFile_32x4__1410_/Q Inst_RegFile_32x4/_0565_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0568_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_my_mux2_inst__1_/A1 ConfigBits\[157\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0964_ Inst_RegFile_32x4__1390_/D Inst_RegFile_32x4__1390_/Q ConfigBits\[1\]
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0417_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0895_ Inst_RegFile_32x4/_0352_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1388_/D
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1447_ net205 Inst_RegFile_32x4/_0099_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1447_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1378_ net205 Inst_RegFile_32x4/_0038_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1378_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix__17_ JN2BEG\[1\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2 BD0 BD1
+ BD2 BD3 ConfigBits\[54\] ConfigBits\[55\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0680_ Inst_RegFile_32x4/_0136_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0146_
+ sky130_fd_sc_hd__buf_2
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1301_ Inst_RegFile_32x4/_0640_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0110_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2 net245
+ AD0 AD1 AD2 ConfigBits\[374\] ConfigBits\[375\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1232_ Inst_RegFile_32x4/_0577_ Inst_RegFile_32x4__1428_/Q Inst_RegFile_32x4/_0601_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XNN4BEG_outbuf_6__0_ NN4BEG_i\[6\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1094_ Inst_RegFile_32x4/_0517_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0026_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1163_ Inst_RegFile_32x4/_0558_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0054_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0947_ Inst_RegFile_32x4__1458_/Q Inst_RegFile_32x4__1454_/Q Inst_RegFile_32x4/_0314_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0878_ Inst_RegFile_32x4__1440_/Q Inst_RegFile_32x4__1436_/Q Inst_RegFile_32x4/_0335_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput391 net391 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput380 net380 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__clkbuf_4
XSS4BEG_outbuf_9__0_ SS4BEG_i\[9\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame3_bit6 net77 net94 VGND VGND VPWR VPWR ConfigBits\[292\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0801_ Inst_RegFile_32x4/_0188_ Inst_RegFile_32x4/_0263_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0264_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0663_ Inst_RegFile_32x4/_0128_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0129_
+ sky130_fd_sc_hd__buf_1
XFILLER_0_43_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0732_ Inst_RegFile_32x4/_0173_ Inst_RegFile_32x4/_0196_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0197_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__1215_ Inst_RegFile_32x4/_0584_ Inst_RegFile_32x4__1423_/Q Inst_RegFile_32x4/_0586_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0590_ sky130_fd_sc_hd__mux2_1
Xinput108 N2END[3] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1077_ Inst_RegFile_32x4/_0507_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0019_
+ sky130_fd_sc_hd__clkbuf_1
Xinput119 N2MID[6] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1146_ Inst_RegFile_32x4/_0548_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0047_
+ sky130_fd_sc_hd__clkbuf_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst1 BD0 J2MID_EFa_BEG\[2\]
+ J2MID_GHa_BEG\[2\] J2END_AB_BEG\[3\] ConfigBits\[83\] ConfigBits\[84\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XNN4END_inbuf_3__0_ net150 VGND VGND VPWR VPWR NN4BEG_i\[3\] sky130_fd_sc_hd__buf_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2 net208
+ AD0 AD1 AD2 ConfigBits\[338\] ConfigBits\[339\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1000_ D0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0450_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0715_ Inst_RegFile_32x4/_0167_ Inst_RegFile_32x4/_0172_ Inst_RegFile_32x4/_0176_
+ Inst_RegFile_32x4/_0180_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0181_ sky130_fd_sc_hd__o22a_1
Xinput90 FrameStrobe[18] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1129_ Inst_RegFile_32x4/_0485_ Inst_RegFile_32x4/_0502_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0539_ sky130_fd_sc_hd__nor2_2
XInst_RegFile_ConfigMem_Inst_frame0_bit9 net80 net81 VGND VGND VPWR VPWR ConfigBits\[391\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3/X ConfigBits\[264\]
+ ConfigBits\[265\] VGND VGND VPWR VPWR JN2BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame9_bit1 net60 net100 VGND VGND VPWR VPWR ConfigBits\[95\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit5 net76 net82 VGND VGND VPWR VPWR ConfigBits\[67\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__50_ JW2BEG\[2\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_1
XN4BEG_outbuf_10__0_ N4BEG_i\[10\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3 AD3 BD1
+ BD2 BD3 ConfigBits\[302\] ConfigBits\[303\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__buf_1
XS4END_inbuf_8__0_ net176 VGND VGND VPWR VPWR S4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0980_ Inst_RegFile_32x4/_0428_ Inst_RegFile_32x4/_0430_ Inst_RegFile_32x4/_0431_
+ Inst_RegFile_32x4/_0310_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0432_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1394_ net205 Inst_RegFile_32x4/_0046_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1394_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1463_ net205 Inst_RegFile_32x4/_0115_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1463_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__33_ JS2BEG\[1\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XEE4BEG_outbuf_9__0_ EE4BEG_i\[9\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame6_bit4 net75 net97 VGND VGND VPWR VPWR ConfigBits\[194\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0963_ Inst_RegFile_32x4/_0416_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1390_/D
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0894_ Inst_RegFile_32x4/_0312_ Inst_RegFile_32x4/_0325_ Inst_RegFile_32x4/_0342_
+ Inst_RegFile_32x4/_0351_ B_ADR3 B_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0352_
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1446_ net205 Inst_RegFile_32x4/_0098_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1446_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1377_ net205 Inst_RegFile_32x4/_0037_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1377_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__16_ JN2BEG\[0\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3 J2MID_ABa_BEG\[2\]
+ J2MID_CDa_BEG\[2\] J2MID_EFa_BEG\[2\] J2MID_GHa_BEG\[2\] ConfigBits\[54\] ConfigBits\[55\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG0 net112 net12 net164 net238
+ ConfigBits\[246\] ConfigBits\[247\] VGND VGND VPWR VPWR J2END_GH_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__1_/A1 ConfigBits\[20\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1300_ Inst_RegFile_32x4__1458_/Q Inst_RegFile_32x4/_0464_ Inst_RegFile_32x4/_0637_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0640_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3 AD3 BD0
+ BD1 BD3 ConfigBits\[374\] ConfigBits\[375\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1231_ Inst_RegFile_32x4/_0570_ Inst_RegFile_32x4/_0600_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0601_ sky130_fd_sc_hd__nand2_2
XInst_RegFile_32x4__1162_ Inst_RegFile_32x4/_0465_ Inst_RegFile_32x4__1402_/Q Inst_RegFile_32x4/_0555_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0558_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1093_ Inst_RegFile_32x4__1366_/Q Inst_RegFile_32x4/_0498_ Inst_RegFile_32x4/_0514_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0517_ sky130_fd_sc_hd__mux2_1
Xdata_inbuf_10__0_ net50 VGND VGND VPWR VPWR FrameData_O_i\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0946_ Inst_RegFile_32x4/_0396_ Inst_RegFile_32x4/_0398_ Inst_RegFile_32x4/_0399_
+ Inst_RegFile_32x4/_0310_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0400_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0877_ Inst_RegFile_32x4/_0291_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0335_
+ sky130_fd_sc_hd__clkbuf_2
Xoutput392 net392 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput381 net381 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput370 net370 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1429_ net205 Inst_RegFile_32x4/_0081_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1429_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame3_bit7 net78 net94 VGND VGND VPWR VPWR ConfigBits\[293\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0731_ Inst_RegFile_32x4__1377_/Q Inst_RegFile_32x4__1373_/Q Inst_RegFile_32x4/_0142_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0196_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0800_ Inst_RegFile_32x4__1363_/Q Inst_RegFile_32x4__1399_/Q Inst_RegFile_32x4/_0136_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0662_ A_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0128_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_28_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1214_ Inst_RegFile_32x4/_0589_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0074_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput109 N2END[4] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1145_ Inst_RegFile_32x4/_0468_ Inst_RegFile_32x4__1395_/Q Inst_RegFile_32x4/_0544_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0548_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1076_ Inst_RegFile_32x4__1359_/Q Inst_RegFile_32x4/_0500_ Inst_RegFile_32x4/_0503_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0507_ sky130_fd_sc_hd__mux2_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0929_ Inst_RegFile_32x4/_0384_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1389_/D
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_60 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_13__0_ FrameStrobe_O_i\[13\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_8__0_ FrameData_O_i\[8\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3 AD3 BD0
+ BD2 BD3 ConfigBits\[338\] ConfigBits\[339\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0714_ Inst_RegFile_32x4/_0145_ Inst_RegFile_32x4/_0178_ Inst_RegFile_32x4/_0179_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0180_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput80 FrameData[9] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_4
Xinput91 FrameStrobe[19] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1128_ Inst_RegFile_32x4/_0538_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0039_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1059_ Inst_RegFile_32x4/_0461_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0496_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XWW4END_inbuf_4__0_ net252 VGND VGND VPWR VPWR WW4BEG_i\[4\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame9_bit2 net71 net100 VGND VGND VPWR VPWR ConfigBits\[96\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit6 net77 net82 VGND VGND VPWR VPWR ConfigBits\[68\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3/X ConfigBits\[304\]
+ ConfigBits\[305\] VGND VGND VPWR VPWR JE2BEG\[4\] sky130_fd_sc_hd__mux4_2
XFILLER_0_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__1_/A1 ConfigBits\[99\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1462_ net205 Inst_RegFile_32x4/_0114_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1462_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1393_ net205 Inst_RegFile_32x4/_0045_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1393_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__32_ JS2BEG\[0\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0 net101
+ net107 net7 net21 ConfigBits\[354\] ConfigBits\[355\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_10__0_ net82 VGND VGND VPWR VPWR FrameStrobe_O_i\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XE6END_inbuf_4__0_ net29 VGND VGND VPWR VPWR E6BEG_i\[4\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame6_bit5 net76 net97 VGND VGND VPWR VPWR ConfigBits\[195\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0893_ Inst_RegFile_32x4/_0345_ Inst_RegFile_32x4/_0348_ Inst_RegFile_32x4/_0350_
+ Inst_RegFile_32x4/_0324_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0351_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_32x4__0962_ Inst_RegFile_32x4/_0394_ Inst_RegFile_32x4/_0400_ Inst_RegFile_32x4/_0409_
+ Inst_RegFile_32x4/_0415_ B_ADR3 B_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0416_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1445_ net205 Inst_RegFile_32x4/_0097_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1445_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__15_ net20 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__1376_ net205 Inst_RegFile_32x4/_0036_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1376_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3/X ConfigBits\[56\]
+ ConfigBits\[57\] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__mux4_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG1 net108 net8 net189 net213
+ ConfigBits\[248\] ConfigBits\[249\] VGND VGND VPWR VPWR J2END_GH_BEG\[1\] sky130_fd_sc_hd__mux4_2
XSS4END_inbuf_6__0_ net190 VGND VGND VPWR VPWR SS4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3/X ConfigBits\[376\]
+ ConfigBits\[377\] VGND VGND VPWR VPWR JW2BEG\[6\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__1230_ W_ADR3 W_ADR2 W_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0600_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1161_ Inst_RegFile_32x4/_0557_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0053_
+ sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_8__0_ FrameStrobe_O_i\[8\] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_1
Xinput1 E1END[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
XInst_RegFile_32x4__1092_ Inst_RegFile_32x4/_0516_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0025_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0876_ Inst_RegFile_32x4/_0289_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0334_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_19_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0945_ Inst_RegFile_32x4__1346_/Q Inst_RegFile_32x4__1394_/Q Inst_RegFile_32x4__1466_/Q
+ Inst_RegFile_32x4__1462_/Q Inst_RegFile_32x4/_0307_ Inst_RegFile_32x4/_0322_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0399_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1428_ net205 Inst_RegFile_32x4/_0080_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1428_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput393 net393 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput382 net382 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput371 net371 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput360 net360 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1359_ net205 Inst_RegFile_32x4/_0019_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1359_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0 net106
+ net4 net6 net24 ConfigBits\[318\] ConfigBits\[319\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame3_bit8 net79 net94 VGND VGND VPWR VPWR ConfigBits\[294\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XEE4END_inbuf_5__0_ net48 VGND VGND VPWR VPWR EE4BEG_i\[5\] sky130_fd_sc_hd__clkbuf_2
Xdata_inbuf_2__0_ net71 VGND VGND VPWR VPWR FrameData_O_i\[2\] sky130_fd_sc_hd__buf_1
XFILLER_0_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XWW4BEG_outbuf_6__0_ WW4BEG_i\[6\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0730_ Inst_RegFile_32x4/_0135_ Inst_RegFile_32x4/_0194_ Inst_RegFile_32x4/_0139_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0195_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_cus_mux41_buf_inst0 net105 net157
+ J2MID_EFa_BEG\[1\] J2MID_EFb_BEG\[2\] ConfigBits\[152\] ConfigBits\[153\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1213_ Inst_RegFile_32x4/_0582_ Inst_RegFile_32x4__1422_/Q Inst_RegFile_32x4/_0586_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1075_ Inst_RegFile_32x4/_0506_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0018_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1144_ Inst_RegFile_32x4/_0547_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0046_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_50 N4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_61 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0859_ Inst_RegFile_32x4/_0291_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0317_
+ sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__0928_ Inst_RegFile_32x4/_0362_ Inst_RegFile_32x4/_0368_ Inst_RegFile_32x4/_0377_
+ Inst_RegFile_32x4/_0383_ B_ADR3 B_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0384_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XE6BEG_outbuf_9__0_ E6BEG_i\[9\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3/X ConfigBits\[340\]
+ ConfigBits\[341\] VGND VGND VPWR VPWR JS2BEG\[5\] sky130_fd_sc_hd__mux4_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0713_ Inst_RegFile_32x4/_0148_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0179_
+ sky130_fd_sc_hd__dlymetal6s2s_1
Xinput70 FrameData[29] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_6
Xinput92 FrameStrobe[1] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_12
XN4END_inbuf_8__0_ net124 VGND VGND VPWR VPWR N4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_2
Xinput81 FrameStrobe[0] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_12
XInst_RegFile_32x4__1127_ Inst_RegFile_32x4__1379_/Q Inst_RegFile_32x4/_0532_ Inst_RegFile_32x4/_0534_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0538_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1058_ Inst_RegFile_32x4/_0495_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0012_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame9_bit3 net74 net100 VGND VGND VPWR VPWR ConfigBits\[97\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit7 net78 net82 VGND VGND VPWR VPWR ConfigBits\[69\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XN4BEG_outbuf_0__0_ N4BEG_i\[0\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst0 net103
+ net155 net208 AD1 ConfigBits\[94\] ConfigBits\[95\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XW6BEG_outbuf_0__0_ W6BEG_i\[0\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1461_ net205 Inst_RegFile_32x4/_0113_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1461_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix__31_ net120 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1392_ net205 Inst_RegFile_32x4/_0044_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1392_/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1 net159
+ net181 net196 net212 ConfigBits\[354\] ConfigBits\[355\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame6_bit6 net77 net97 VGND VGND VPWR VPWR ConfigBits\[196\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0961_ Inst_RegFile_32x4/_0411_ Inst_RegFile_32x4/_0413_ Inst_RegFile_32x4/_0414_
+ Inst_RegFile_32x4/_0324_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0415_ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0892_ Inst_RegFile_32x4__1408_/Q Inst_RegFile_32x4__1340_/Q Inst_RegFile_32x4__1400_/Q
+ Inst_RegFile_32x4__1468_/Q Inst_RegFile_32x4/_0321_ Inst_RegFile_32x4/_0349_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0350_ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1444_ net205 Inst_RegFile_32x4/_0096_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1444_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XNN4BEG_outbuf_9__0_ NN4BEG_i\[9\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_outbuf_20__0_ FrameData_O_i\[20\] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix__14_ net19 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__1375_ net205 Inst_RegFile_32x4/_0035_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1375_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG2 net144 net10 net162 net215
+ ConfigBits\[250\] ConfigBits\[251\] VGND VGND VPWR VPWR J2END_GH_BEG\[2\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0 net109
+ net121 net3 net9 ConfigBits\[266\] ConfigBits\[267\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_outbuf_11__0_ FrameData_O_i\[11\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XS4BEG_outbuf_0__0_ S4BEG_i\[0\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1091_ Inst_RegFile_32x4__1365_/Q Inst_RegFile_32x4/_0496_ Inst_RegFile_32x4/_0514_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1160_ Inst_RegFile_32x4/_0462_ Inst_RegFile_32x4__1401_/Q Inst_RegFile_32x4/_0555_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0557_ sky130_fd_sc_hd__mux2_1
Xinput2 E1END[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0875_ Inst_RegFile_32x4/_0329_ Inst_RegFile_32x4/_0331_ Inst_RegFile_32x4/_0332_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0333_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0944_ Inst_RegFile_32x4/_0302_ Inst_RegFile_32x4/_0397_ Inst_RegFile_32x4/_0319_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0398_ sky130_fd_sc_hd__a21o_1
Xoutput350 net350 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__clkbuf_4
Xoutput361 net361 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1427_ net205 Inst_RegFile_32x4/_0079_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1427_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1358_ net205 Inst_RegFile_32x4/_0018_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1358_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput372 net372 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput394 net394 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput383 net383 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1289_ Inst_RegFile_32x4__1453_/Q Inst_RegFile_32x4/_0594_ Inst_RegFile_32x4/_0632_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0634_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1 net158
+ net180 net211 net238 ConfigBits\[318\] ConfigBits\[319\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame3_bit9 net80 net94 VGND VGND VPWR VPWR ConfigBits\[295\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_cus_mux41_buf_inst1 J2END_AB_BEG\[3\]
+ JN2BEG\[7\] JS2BEG\[7\] JW2BEG\[7\] ConfigBits\[152\] ConfigBits\[153\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1212_ Inst_RegFile_32x4/_0588_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0073_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XNN4END_inbuf_6__0_ net138 VGND VGND VPWR VPWR NN4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1074_ Inst_RegFile_32x4__1358_/Q Inst_RegFile_32x4/_0498_ Inst_RegFile_32x4/_0503_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XW6END_inbuf_2__0_ net232 VGND VGND VPWR VPWR W6BEG_i\[2\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1143_ Inst_RegFile_32x4/_0465_ Inst_RegFile_32x4__1394_/Q Inst_RegFile_32x4/_0544_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0547_ sky130_fd_sc_hd__mux2_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0927_ Inst_RegFile_32x4/_0379_ Inst_RegFile_32x4/_0381_ Inst_RegFile_32x4/_0382_
+ Inst_RegFile_32x4/_0324_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0383_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_62 JN2BEG\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 NN4BEG_i\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG0 net111 net11 net198 net216
+ ConfigBits\[222\] ConfigBits\[223\] VGND VGND VPWR VPWR J2END_AB_BEG\[0\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0789_ Inst_RegFile_32x4/_0231_ Inst_RegFile_32x4/_0237_ Inst_RegFile_32x4/_0246_
+ Inst_RegFile_32x4/_0252_ A_ADR3 A_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0253_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_40 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0858_ Inst_RegFile_32x4/_0313_ Inst_RegFile_32x4/_0315_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0316_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst0 net101
+ net1 net153 AD3 ConfigBits\[44\] ConfigBits\[45\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0712_ Inst_RegFile_32x4__1432_/Q Inst_RegFile_32x4__1428_/Q Inst_RegFile_32x4/_0177_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput71 FrameData[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_8
Xinput60 FrameData[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_4
XFILLER_0_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput93 FrameStrobe[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_12
Xinput82 FrameStrobe[10] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_12
XFILLER_0_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1126_ Inst_RegFile_32x4/_0537_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0038_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1057_ Inst_RegFile_32x4__1352_/Q Inst_RegFile_32x4/_0491_ Inst_RegFile_32x4/_0494_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame9_bit4 net75 net100 VGND VGND VPWR VPWR ConfigBits\[98\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit8 net79 net82 VGND VGND VPWR VPWR ConfigBits\[70\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1109_ Inst_RegFile_32x4__1372_/Q Inst_RegFile_32x4/_0524_ Inst_RegFile_32x4/_0526_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput250 WW4END[6] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst1 BD1 J2MID_ABb_BEG\[1\]
+ J2MID_CDb_BEG\[1\] J2END_GH_BEG\[2\] ConfigBits\[94\] ConfigBits\[95\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1391_ net205 Inst_RegFile_32x4__1391_/D VGND VGND VPWR VPWR Inst_RegFile_32x4__1391_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1460_ net205 Inst_RegFile_32x4/_0112_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1460_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix__30_ net119 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2 net226
+ AD0 AD2 AD3 ConfigBits\[354\] ConfigBits\[355\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
Xdata_inbuf_31__0_ net73 VGND VGND VPWR VPWR FrameData_O_i\[31\] sky130_fd_sc_hd__buf_1
XInst_RegFile_ConfigMem_Inst_frame6_bit7 net78 net97 VGND VGND VPWR VPWR ConfigBits\[197\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0960_ Inst_RegFile_32x4__1410_/Q Inst_RegFile_32x4__1342_/Q Inst_RegFile_32x4__1402_/Q
+ Inst_RegFile_32x4__1470_/Q Inst_RegFile_32x4/_0321_ Inst_RegFile_32x4/_0322_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0414_ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_N1BEG0 AD2 J2MID_CDb_BEG\[3\] JW2BEG\[3\]
+ J_l_CD_BEG\[1\] ConfigBits\[2\] ConfigBits\[3\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__mux4_2
XFILLER_0_73_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_22__0_ net63 VGND VGND VPWR VPWR FrameData_O_i\[22\] sky130_fd_sc_hd__buf_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0891_ B_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0349_ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_32x4__1443_ net205 Inst_RegFile_32x4/_0095_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1443_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1374_ net205 Inst_RegFile_32x4/_0034_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1374_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix__13_ net18 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG3 net106 net42 net158 net211
+ ConfigBits\[252\] ConfigBits\[253\] VGND VGND VPWR VPWR J2END_GH_BEG\[3\] sky130_fd_sc_hd__mux4_2
Xstrobe_inbuf_1__0_ net92 VGND VGND VPWR VPWR FrameStrobe_O_i\[1\] sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_13__0_ net53 VGND VGND VPWR VPWR FrameData_O_i\[13\] sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1 net21
+ net161 net214 net247 ConfigBits\[266\] ConfigBits\[267\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XWW4BEG_outbuf_10__0_ WW4BEG_i\[10\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1090_ Inst_RegFile_32x4/_0515_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0024_
+ sky130_fd_sc_hd__clkbuf_1
Xinput3 E1END[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_36_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0943_ Inst_RegFile_32x4__1354_/Q Inst_RegFile_32x4__1350_/Q Inst_RegFile_32x4/_0303_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0397_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0 net103
+ net111 net3 net11 ConfigBits\[306\] ConfigBits\[307\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0874_ B_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0332_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput351 net351 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__clkbuf_4
Xoutput395 net395 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput384 net384 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput373 net373 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput362 net362 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput340 net340 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1426_ net205 Inst_RegFile_32x4/_0078_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1426_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1357_ net205 Inst_RegFile_32x4/_0017_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1357_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2 net229
+ AD1 AD2 AD3 ConfigBits\[318\] ConfigBits\[319\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1288_ Inst_RegFile_32x4/_0633_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0104_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_W_ADR0 J2MID_CDa_BEG\[0\] J2MID_CDb_BEG\[0\]
+ J2END_CD_BEG\[0\] J_l_CD_BEG\[0\] ConfigBits\[144\] ConfigBits\[145\] VGND VGND
+ VPWR VPWR W_ADR0 sky130_fd_sc_hd__mux4_2
Xstrobe_outbuf_16__0_ FrameStrobe_O_i\[16\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1211_ Inst_RegFile_32x4/_0580_ Inst_RegFile_32x4__1421_/Q Inst_RegFile_32x4/_0586_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0588_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1073_ Inst_RegFile_32x4/_0505_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0017_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1142_ Inst_RegFile_32x4/_0546_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0045_
+ sky130_fd_sc_hd__clkbuf_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0926_ Inst_RegFile_32x4__1409_/Q Inst_RegFile_32x4__1341_/Q Inst_RegFile_32x4__1401_/Q
+ Inst_RegFile_32x4__1469_/Q Inst_RegFile_32x4/_0321_ Inst_RegFile_32x4/_0349_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0382_ sky130_fd_sc_hd__mux4_1
XANTENNA_63 NN4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0788_ Inst_RegFile_32x4/_0248_ Inst_RegFile_32x4/_0250_ Inst_RegFile_32x4/_0251_
+ Inst_RegFile_32x4/_0163_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0252_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG1 net137 net7 net159 net212
+ ConfigBits\[224\] ConfigBits\[225\] VGND VGND VPWR VPWR J2END_AB_BEG\[1\] sky130_fd_sc_hd__mux4_2
XANTENNA_41 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0857_ Inst_RegFile_32x4__1360_/Q Inst_RegFile_32x4__1396_/Q Inst_RegFile_32x4/_0314_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0315_ sky130_fd_sc_hd__mux2_1
XANTENNA_52 S4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinst_clk_buf net205 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1409_ net205 Inst_RegFile_32x4/_0061_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1409_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XWW4END_inbuf_7__0_ net240 VGND VGND VPWR VPWR WW4BEG_i\[7\] sky130_fd_sc_hd__clkbuf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst1 BD3 J2MID_EFb_BEG\[1\]
+ J2MID_GHb_BEG\[1\] J2END_CD_BEG\[0\] ConfigBits\[44\] ConfigBits\[45\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0711_ Inst_RegFile_32x4/_0136_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0177_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput72 FrameData[30] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_8
Xinput61 FrameData[20] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput50 FrameData[10] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1125_ Inst_RegFile_32x4__1378_/Q Inst_RegFile_32x4/_0530_ Inst_RegFile_32x4/_0534_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0537_ sky130_fd_sc_hd__mux2_1
Xinput94 FrameStrobe[3] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_16
Xinput83 FrameStrobe[11] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_12
XInst_RegFile_32x4__1056_ Inst_RegFile_32x4/_0483_ Inst_RegFile_32x4/_0493_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0494_ sky130_fd_sc_hd__nor2_2
XInst_RegFile_32x4__0909_ Inst_RegFile_32x4__1353_/Q Inst_RegFile_32x4__1349_/Q Inst_RegFile_32x4/_0317_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0 net101
+ net105 net1 net5 ConfigBits\[378\] ConfigBits\[379\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame9_bit5 net76 net100 VGND VGND VPWR VPWR ConfigBits\[99\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit9 net80 net82 VGND VGND VPWR VPWR ConfigBits\[71\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_53_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1108_ Inst_RegFile_32x4/_0525_ Inst_RegFile_32x4/_0513_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0526_ sky130_fd_sc_hd__nor2_2
XFILLER_0_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG0 net130 net8 net213 JN2BEG\[3\]
+ ConfigBits\[398\] ConfigBits\[399\] VGND VGND VPWR VPWR J_l_EF_BEG\[0\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1039_ Inst_RegFile_32x4__1347_/Q Inst_RegFile_32x4/_0481_ Inst_RegFile_32x4/_0475_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_13__0_ net85 VGND VGND VPWR VPWR FrameStrobe_O_i\[13\] sky130_fd_sc_hd__clkbuf_2
XE6END_inbuf_7__0_ net32 VGND VGND VPWR VPWR E6BEG_i\[7\] sky130_fd_sc_hd__clkbuf_2
Xinput240 WW4END[11] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
Xinput251 WW4END[7] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1390_ net205 Inst_RegFile_32x4__1390_/D VGND VGND VPWR VPWR Inst_RegFile_32x4__1390_/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[354\] ConfigBits\[355\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XSS4END_inbuf_9__0_ net193 VGND VGND VPWR VPWR SS4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0 net104
+ net112 net4 net12 ConfigBits\[342\] ConfigBits\[343\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame6_bit8 net79 net97 VGND VGND VPWR VPWR ConfigBits\[198\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0890_ Inst_RegFile_32x4/_0346_ Inst_RegFile_32x4/_0347_ Inst_RegFile_32x4/_0300_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0348_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_N1BEG1 AD3 J2MID_EFb_BEG\[0\] JW2BEG\[0\]
+ J_l_EF_BEG\[2\] ConfigBits\[4\] ConfigBits\[5\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__mux4_2
XFILLER_0_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1442_ net205 Inst_RegFile_32x4/_0094_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1442_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1373_ net205 Inst_RegFile_32x4/_0033_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1373_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput500 net500 VGND VGND VPWR VPWR WW4BEG[3] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix__12_ net17 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2 net226
+ AD0 AD1 AD2 ConfigBits\[266\] ConfigBits\[267\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XEE4END_inbuf_8__0_ net36 VGND VGND VPWR VPWR EE4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_2
Xdata_inbuf_5__0_ net76 VGND VGND VPWR VPWR FrameData_O_i\[5\] sky130_fd_sc_hd__buf_1
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 E1END[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_8
XWW4BEG_outbuf_9__0_ WW4BEG_i\[9\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0873_ Inst_RegFile_32x4__1448_/Q Inst_RegFile_32x4__1472_/Q Inst_RegFile_32x4/_0330_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0331_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0942_ Inst_RegFile_32x4/_0349_ Inst_RegFile_32x4/_0395_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0396_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1 net41
+ net153 net155 net163 ConfigBits\[306\] ConfigBits\[307\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput352 net352 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__clkbuf_4
Xoutput385 net385 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput396 net396 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput374 net374 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput363 net363 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1287_ Inst_RegFile_32x4__1452_/Q Inst_RegFile_32x4/_0591_ Inst_RegFile_32x4/_0632_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0633_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1425_ net205 Inst_RegFile_32x4/_0077_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1425_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput330 net330 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1356_ net205 Inst_RegFile_32x4/_0016_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1356_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[318\] ConfigBits\[319\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_W_ADR1 J2MID_CDa_BEG\[1\] J2MID_CDb_BEG\[1\]
+ J2END_CD_BEG\[1\] J_l_CD_BEG\[1\] ConfigBits\[146\] ConfigBits\[147\] VGND VGND
+ VPWR VPWR W_ADR1 sky130_fd_sc_hd__mux4_1
XFILLER_0_28_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1210_ Inst_RegFile_32x4/_0587_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0072_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1141_ Inst_RegFile_32x4/_0462_ Inst_RegFile_32x4__1393_/Q Inst_RegFile_32x4/_0544_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0546_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1072_ Inst_RegFile_32x4__1357_/Q Inst_RegFile_32x4/_0496_ Inst_RegFile_32x4/_0503_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_20 NN4BEG_i\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0856_ B_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0314_ sky130_fd_sc_hd__buf_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0925_ Inst_RegFile_32x4/_0346_ Inst_RegFile_32x4/_0380_ Inst_RegFile_32x4/_0332_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0381_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_ConfigMem_Inst_frame2_bit0 net49 net93 VGND VGND VPWR VPWR ConfigBits\[318\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG2 net109 net33 net161 net214
+ ConfigBits\[226\] ConfigBits\[227\] VGND VGND VPWR VPWR J2END_AB_BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_42 net263 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_53 SS4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 S4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0787_ Inst_RegFile_32x4__1410_/Q Inst_RegFile_32x4__1342_/Q Inst_RegFile_32x4__1402_/Q
+ Inst_RegFile_32x4__1470_/Q Inst_RegFile_32x4/_0160_ Inst_RegFile_32x4/_0161_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0251_ sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__1408_ net205 Inst_RegFile_32x4/_0060_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1408_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1339_ Inst_RegFile_32x4/_0661_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0127_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XN4BEG_outbuf_3__0_ N4BEG_i\[3\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0710_ Inst_RegFile_32x4/_0173_ Inst_RegFile_32x4/_0175_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0176_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput73 FrameData[31] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput62 FrameData[21] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_8
Xinput51 FrameData[11] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_6
Xinput40 EE4END[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XFILLER_0_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput95 FrameStrobe[4] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_16
Xinput84 FrameStrobe[12] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_16
XInst_RegFile_32x4__1124_ Inst_RegFile_32x4/_0536_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0037_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1055_ Inst_RegFile_32x4/_0484_ Inst_RegFile_32x4/_0492_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0493_ sky130_fd_sc_hd__or2_2
XSS4BEG_outbuf_2__0_ SS4BEG_i\[2\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0839_ B_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0297_ sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__0908_ Inst_RegFile_32x4/_0349_ Inst_RegFile_32x4/_0363_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0364_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame9_bit6 net77 net100 VGND VGND VPWR VPWR ConfigBits\[100\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XSS4BEG_outbuf_10__0_ SS4BEG_i\[10\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1 net153
+ net155 net157 net206 ConfigBits\[378\] ConfigBits\[379\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XW6BEG_outbuf_3__0_ W6BEG_i\[3\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1107_ Inst_RegFile_32x4/_0456_ Inst_RegFile_32x4/_0484_ Inst_RegFile_32x4/_0457_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0525_ sky130_fd_sc_hd__nand3b_4
XInst_RegFile_32x4__1038_ D3 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0481_ sky130_fd_sc_hd__buf_1
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG1 net145 net7 net181 JE2BEG\[3\]
+ ConfigBits\[400\] ConfigBits\[401\] VGND VGND VPWR VPWR J_l_EF_BEG\[1\] sky130_fd_sc_hd__mux4_1
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput230 W6END[2] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
Xinput241 WW4END[12] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_1
Xinput252 WW4END[8] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_outbuf_23__0_ FrameData_O_i\[23\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3/X ConfigBits\[356\]
+ ConfigBits\[357\] VGND VGND VPWR VPWR JW2BEG\[1\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame6_bit9 net80 net97 VGND VGND VPWR VPWR ConfigBits\[199\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1 net156
+ net164 net196 net207 ConfigBits\[342\] ConfigBits\[343\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_outbuf_14__0_ FrameData_O_i\[14\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_N1BEG2 BD0 J2MID_GHb_BEG\[1\] JW2BEG\[1\]
+ J_l_GH_BEG\[3\] ConfigBits\[6\] ConfigBits\[7\] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__mux4_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4BEG_outbuf_3__0_ S4BEG_i\[3\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1441_ net205 Inst_RegFile_32x4/_0093_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1441_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix__11_ net16 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1372_ net205 Inst_RegFile_32x4/_0032_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1372_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput501 net501 VGND VGND VPWR VPWR WW4BEG[4] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[266\] ConfigBits\[267\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XS4END_inbuf_1__0_ net184 VGND VGND VPWR VPWR S4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput5 E2END[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0872_ Inst_RegFile_32x4/_0291_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0330_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0941_ Inst_RegFile_32x4__1362_/Q Inst_RegFile_32x4__1398_/Q Inst_RegFile_32x4/_0314_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0395_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2 net208
+ AD0 AD1 AD2 ConfigBits\[306\] ConfigBits\[307\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1424_ net205 Inst_RegFile_32x4/_0076_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1424_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XNN4END_inbuf_9__0_ net141 VGND VGND VPWR VPWR NN4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput364 net364 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput353 net353 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput397 net397 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput386 net386 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput375 net375 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput320 net320 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput331 net331 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__clkbuf_4
XEE4BEG_outbuf_2__0_ EE4BEG_i\[2\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1286_ Inst_RegFile_32x4/_0525_ Inst_RegFile_32x4/_0626_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0632_ sky130_fd_sc_hd__nor2_2
XW6END_inbuf_5__0_ net235 VGND VGND VPWR VPWR W6BEG_i\[5\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3/X ConfigBits\[320\]
+ ConfigBits\[321\] VGND VGND VPWR VPWR JS2BEG\[0\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__1355_ net205 Inst_RegFile_32x4/_0015_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1355_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG0 net120 net20 net172
+ net225 ConfigBits\[206\] ConfigBits\[207\] VGND VGND VPWR VPWR J2MID_EFb_BEG\[0\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame12_bit30 net72 net84 VGND VGND VPWR VPWR ConfigBits\[28\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_W_ADR2 J2MID_CDa_BEG\[2\] J2MID_CDb_BEG\[2\]
+ J2END_CD_BEG\[2\] J_l_CD_BEG\[2\] ConfigBits\[148\] ConfigBits\[149\] VGND VGND
+ VPWR VPWR W_ADR2 sky130_fd_sc_hd__mux4_2
XFILLER_0_24_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1071_ Inst_RegFile_32x4/_0504_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0016_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1140_ Inst_RegFile_32x4/_0545_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0044_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_32 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 E6BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0786_ Inst_RegFile_32x4/_0185_ Inst_RegFile_32x4/_0249_ Inst_RegFile_32x4/_0171_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0250_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0924_ Inst_RegFile_32x4__1417_/Q Inst_RegFile_32x4__1413_/Q Inst_RegFile_32x4/_0330_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0380_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG3 net105 net5 net157 net247
+ ConfigBits\[228\] ConfigBits\[229\] VGND VGND VPWR VPWR J2END_AB_BEG\[3\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__0855_ Inst_RegFile_32x4/_0289_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0313_
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_54 SS4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 S4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_ConfigMem_Inst_frame2_bit1 net60 net93 VGND VGND VPWR VPWR ConfigBits\[319\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_10 JW2BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1407_ net205 Inst_RegFile_32x4/_0059_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1407_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1338_ Inst_RegFile_32x4__1475_/Q Inst_RegFile_32x4/_0467_ Inst_RegFile_32x4/_0657_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0661_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1269_ Inst_RegFile_32x4/_0622_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0096_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput63 FrameData[22] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_8
Xinput52 FrameData[12] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_8
Xinput74 FrameData[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_8
Xinput30 E6END[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 EE4END[2] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput96 FrameStrobe[5] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_16
Xinput85 FrameStrobe[13] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1123_ Inst_RegFile_32x4__1377_/Q Inst_RegFile_32x4/_0528_ Inst_RegFile_32x4/_0534_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0536_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1054_ Inst_RegFile_32x4/_0456_ Inst_RegFile_32x4/_0457_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0907_ Inst_RegFile_32x4__1361_/Q Inst_RegFile_32x4__1397_/Q Inst_RegFile_32x4/_0314_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0363_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0838_ Inst_RegFile_32x4/_0295_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0296_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0769_ Inst_RegFile_32x4/_0188_ Inst_RegFile_32x4/_0232_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0233_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2 net238
+ AD0 AD1 AD2 ConfigBits\[378\] ConfigBits\[379\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame9_bit7 net78 net100 VGND VGND VPWR VPWR ConfigBits\[101\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1106_ D0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0524_ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_32x4__1037_ Inst_RegFile_32x4/_0480_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0006_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG2 net128 net196 net214 JS2BEG\[3\]
+ ConfigBits\[402\] ConfigBits\[403\] VGND VGND VPWR VPWR J_l_EF_BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_1__0_ FrameData_O_i\[1\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_1
Xinput231 W6END[3] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_1
Xinput242 WW4END[13] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_1
Xinput253 WW4END[9] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_1
Xinput220 W2MID[2] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_inbuf_25__0_ net66 VGND VGND VPWR VPWR FrameData_O_i\[25\] sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_N4BEG0 net107 net128 net24 BD0 ConfigBits\[10\]
+ ConfigBits\[11\] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__mux4_2
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_4__0_ net95 VGND VGND VPWR VPWR FrameStrobe_O_i\[4\] sky130_fd_sc_hd__clkbuf_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_inbuf_16__0_ net56 VGND VGND VPWR VPWR FrameData_O_i\[16\] sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2 net209
+ AD0 AD1 AD2 ConfigBits\[342\] ConfigBits\[343\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_N1BEG3 BD1 J2MID_ABb_BEG\[2\] JW2BEG\[2\]
+ J_l_AB_BEG\[0\] ConfigBits\[8\] ConfigBits\[9\] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__mux4_1
XFILLER_0_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1440_ net205 Inst_RegFile_32x4/_0092_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1440_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1371_ net205 Inst_RegFile_32x4/_0031_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1371_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput502 net502 VGND VGND VPWR VPWR WW4BEG[5] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix__10_ net15 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__buf_1
XFILLER_0_22_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3/X ConfigBits\[268\]
+ ConfigBits\[269\] VGND VGND VPWR VPWR JN2BEG\[3\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG0 net19 net171 net224
+ JN2BEG\[4\] ConfigBits\[166\] ConfigBits\[167\] VGND VGND VPWR VPWR J2MID_CDa_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xstrobe_outbuf_19__0_ FrameStrobe_O_i\[19\] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0940_ Inst_RegFile_32x4/_0387_ Inst_RegFile_32x4/_0389_ Inst_RegFile_32x4/_0391_
+ Inst_RegFile_32x4/_0393_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0394_ sky130_fd_sc_hd__o22a_1
Xinput6 E2END[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0871_ Inst_RegFile_32x4/_0295_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0329_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput343 net343 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput321 net321 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3 AD3 BD0
+ BD2 BD3 ConfigBits\[306\] ConfigBits\[307\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xoutput310 net310 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput332 net332 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1423_ net205 Inst_RegFile_32x4/_0075_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1423_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1354_ net205 Inst_RegFile_32x4/_0014_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1354_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput387 net387 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput398 net398 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput376 net376 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput365 net365 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1285_ Inst_RegFile_32x4/_0631_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0103_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG1 net116 net16 net168
+ net221 ConfigBits\[208\] ConfigBits\[209\] VGND VGND VPWR VPWR J2MID_EFb_BEG\[1\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame12_bit20 net61 net84 VGND VGND VPWR VPWR ConfigBits\[18\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit31 net73 net84 VGND VGND VPWR VPWR ConfigBits\[29\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_W_ADR3 J2MID_CDa_BEG\[3\] J2MID_CDb_BEG\[3\]
+ J2END_CD_BEG\[3\] J_l_CD_BEG\[3\] ConfigBits\[150\] ConfigBits\[151\] VGND VGND
+ VPWR VPWR W_ADR3 sky130_fd_sc_hd__mux4_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1070_ Inst_RegFile_32x4__1356_/Q Inst_RegFile_32x4/_0491_ Inst_RegFile_32x4/_0503_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0504_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0923_ Inst_RegFile_32x4/_0343_ ANTENNA_55/DIODE VGND VGND VPWR
+ VPWR Inst_RegFile_32x4/_0379_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_44 J2MID_EFb_BEG\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0785_ Inst_RegFile_32x4__1418_/Q Inst_RegFile_32x4__1414_/Q Inst_RegFile_32x4/_0169_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0249_ sky130_fd_sc_hd__mux2_1
XANTENNA_55 ANTENNA_55/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0854_ Inst_RegFile_32x4/_0294_ Inst_RegFile_32x4/_0301_ Inst_RegFile_32x4/_0305_
+ Inst_RegFile_32x4/_0311_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0312_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_22 S4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_ConfigMem_Inst_frame2_bit2 net71 net93 VGND VGND VPWR VPWR ConfigBits\[320\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_11 JW2BEG\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__1337_ Inst_RegFile_32x4/_0660_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0126_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1406_ net205 Inst_RegFile_32x4/_0058_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1406_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1199_ Inst_RegFile_32x4/_0461_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0580_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_32x4__1268_ Inst_RegFile_32x4__1444_/Q Inst_RegFile_32x4/_0591_ Inst_RegFile_32x4/_0621_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_1__0_ FrameStrobe_O_i\[1\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput31 E6END[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 E2MID[7] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
Xinput64 FrameData[23] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_8
Xinput53 FrameData[13] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_8
Xinput75 FrameData[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_8
Xinput42 EE4END[3] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput97 FrameStrobe[6] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_16
Xinput86 FrameStrobe[14] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1053_ Inst_RegFile_32x4/_0450_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0491_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1122_ Inst_RegFile_32x4/_0535_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0036_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0906_ Inst_RegFile_32x4/_0355_ Inst_RegFile_32x4/_0357_ Inst_RegFile_32x4/_0359_
+ Inst_RegFile_32x4/_0361_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0362_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0699_ A_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0165_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame11_bit30 net72 net83 VGND VGND VPWR VPWR ConfigBits\[60\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0837_ B_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0295_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0768_ Inst_RegFile_32x4__1362_/Q Inst_RegFile_32x4__1398_/Q Inst_RegFile_32x4/_0153_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0232_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3 AD3 BD0
+ BD1 BD2 ConfigBits\[378\] ConfigBits\[379\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame9_bit8 net79 net100 VGND VGND VPWR VPWR ConfigBits\[102\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xstrobe_inbuf_16__0_ net88 VGND VGND VPWR VPWR FrameStrobe_O_i\[16\] sky130_fd_sc_hd__clkbuf_2
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1105_ Inst_RegFile_32x4/_0523_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0031_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1036_ Inst_RegFile_32x4__1346_/Q Inst_RegFile_32x4/_0479_ Inst_RegFile_32x4/_0475_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG3 net42 net173 net245 JW2BEG\[3\]
+ ConfigBits\[404\] ConfigBits\[405\] VGND VGND VPWR VPWR J_l_EF_BEG\[3\] sky130_fd_sc_hd__mux4_1
XE6BEG_outbuf_2__0_ E6BEG_i\[2\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_1
Xinput232 W6END[4] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
Xinput243 WW4END[14] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_1
Xinput221 W2MID[3] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_4
Xinput210 W2END[0] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_N4BEG1 net108 net129 net21 BD1 ConfigBits\[12\]
+ ConfigBits\[13\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__mux4_1
XN4END_inbuf_1__0_ net132 VGND VGND VPWR VPWR N4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_2
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1019_ Inst_RegFile_32x4/_0466_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0002_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3 AD3 BD0
+ BD1 BD3 ConfigBits\[342\] ConfigBits\[343\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0 net104
+ net106 net128 net137 ConfigBits\[286\] ConfigBits\[287\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_8__0_ net79 VGND VGND VPWR VPWR FrameData_O_i\[8\] sky130_fd_sc_hd__buf_1
XFILLER_0_58_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1370_ net205 Inst_RegFile_32x4/_0030_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1370_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput503 net503 VGND VGND VPWR VPWR WW4BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__1_/A1 ConfigBits\[46\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame5_bit0 net49 net96 VGND VGND VPWR VPWR ConfigBits\[222\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG1 net115 net15 net220
+ JE2BEG\[4\] ConfigBits\[168\] ConfigBits\[169\] VGND VGND VPWR VPWR J2MID_CDa_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 E2END[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3/X ConfigBits\[308\]
+ ConfigBits\[309\] VGND VGND VPWR VPWR JE2BEG\[5\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__0870_ Inst_RegFile_32x4/_0313_ Inst_RegFile_32x4/_0327_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0328_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput377 net377 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput366 net366 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput355 net355 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput344 net344 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput322 net322 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1284_ Inst_RegFile_32x4__1451_/Q Inst_RegFile_32x4/_0598_ Inst_RegFile_32x4/_0627_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0631_ sky130_fd_sc_hd__mux2_1
Xoutput311 net311 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput333 net333 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1422_ net205 Inst_RegFile_32x4/_0074_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1422_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput300 net300 VGND VGND VPWR VPWR EE4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1353_ net205 Inst_RegFile_32x4/_0013_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1353_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput399 net399 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput388 net388 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG2 net118 net18 net170
+ net223 ConfigBits\[210\] ConfigBits\[211\] VGND VGND VPWR VPWR J2MID_EFb_BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0999_ Inst_RegFile_32x4/_0449_ VGND VGND VPWR VPWR BD3 sky130_fd_sc_hd__buf_12
XFILLER_0_33_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame12_bit21 net62 net84 VGND VGND VPWR VPWR ConfigBits\[19\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit10 net50 net84 VGND VGND VPWR VPWR ConfigBits\[8\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XNN4BEG_outbuf_2__0_ NN4BEG_i\[2\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0 net102
+ net108 net145 net8 ConfigBits\[358\] ConfigBits\[359\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XN4BEG_outbuf_6__0_ N4BEG_i\[6\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0922_ Inst_RegFile_32x4__1425_/Q Inst_RegFile_32x4__1421_/Q Inst_RegFile_32x4/_0326_
+ VGND VGND VPWR VPWR ANTENNA_55/DIODE sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0853_ Inst_RegFile_32x4/_0306_ Inst_RegFile_32x4/_0308_ Inst_RegFile_32x4/_0310_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0311_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_ConfigMem_Inst_frame2_bit3 net74 net93 VGND VGND VPWR VPWR ConfigBits\[321\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0784_ Inst_RegFile_32x4/_0182_ Inst_RegFile_32x4/_0247_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0248_ sky130_fd_sc_hd__and2b_1
XANTENNA_12 JW2BEG\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 JN2BEG\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_23 S4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_34 net146 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__1336_ Inst_RegFile_32x4__1474_/Q Inst_RegFile_32x4/_0464_ Inst_RegFile_32x4/_0657_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0660_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1267_ Inst_RegFile_32x4/_0525_ Inst_RegFile_32x4/_0502_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0621_ sky130_fd_sc_hd__nor2_2
XInst_RegFile_32x4__1405_ net205 Inst_RegFile_32x4/_0057_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1405_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSS4BEG_outbuf_5__0_ SS4BEG_i\[5\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1198_ Inst_RegFile_32x4/_0579_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0068_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput54 FrameData[14] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 E6END[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput21 E6END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput43 EE4END[4] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput10 E2END[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput65 FrameData[24] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_8
Xinput76 FrameData[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_6
XInst_RegFile_32x4__1121_ Inst_RegFile_32x4__1376_/Q Inst_RegFile_32x4/_0524_ Inst_RegFile_32x4/_0534_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0535_ sky130_fd_sc_hd__mux2_1
Xinput98 FrameStrobe[7] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_8
Xinput87 FrameStrobe[15] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XW6BEG_outbuf_6__0_ W6BEG_i\[6\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1052_ Inst_RegFile_32x4/_0490_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0011_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0836_ Inst_RegFile_32x4/_0290_ Inst_RegFile_32x4/_0293_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0294_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0905_ Inst_RegFile_32x4/_0306_ Inst_RegFile_32x4/_0360_ Inst_RegFile_32x4/_0310_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0361_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_ConfigMem_Inst_frame11_bit20 net61 net83 VGND VGND VPWR VPWR ConfigBits\[50\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0767_ Inst_RegFile_32x4/_0224_ Inst_RegFile_32x4/_0226_ Inst_RegFile_32x4/_0228_
+ Inst_RegFile_32x4/_0230_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0231_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_32x4__0698_ Inst_RegFile_32x4/_0155_ Inst_RegFile_32x4/_0159_ Inst_RegFile_32x4/_0162_
+ Inst_RegFile_32x4/_0163_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0164_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_ConfigMem_Inst_frame11_bit31 net73 net83 VGND VGND VPWR VPWR ConfigBits\[61\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1319_ Inst_RegFile_32x4/_0650_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0118_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3/X ConfigBits\[380\]
+ ConfigBits\[381\] VGND VGND VPWR VPWR JW2BEG\[7\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame9_bit9 net80 net100 VGND VGND VPWR VPWR ConfigBits\[103\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__1_/A1 ConfigBits\[29\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0 net107
+ net1 net7 net21 ConfigBits\[322\] ConfigBits\[323\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1104_ Inst_RegFile_32x4__1371_/Q Inst_RegFile_32x4/_0500_ Inst_RegFile_32x4/_0519_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1035_ D2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0479_ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_32x4__0819_ Inst_RegFile_32x4__1411_/Q Inst_RegFile_32x4__1343_/Q Inst_RegFile_32x4__1403_/Q
+ Inst_RegFile_32x4__1471_/Q Inst_RegFile_32x4/_0160_ Inst_RegFile_32x4/_0161_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0282_ sky130_fd_sc_hd__mux4_2
Xdata_outbuf_26__0_ FrameData_O_i\[26\] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__buf_1
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput200 SS4END[5] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
Xinput233 W6END[5] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
Xinput244 WW4END[15] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
Xinput222 W2MID[4] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_2
Xinput211 W2END[1] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_2
XFILLER_0_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_17__0_ FrameData_O_i\[17\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_N4BEG2 net105 net130 net229 BD2 ConfigBits\[14\]
+ ConfigBits\[15\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__mux4_1
XFILLER_0_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XS4BEG_outbuf_6__0_ S4BEG_i\[6\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame10_bit30 net72 net82 VGND VGND VPWR VPWR ConfigBits\[92\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1018_ Inst_RegFile_32x4/_0465_ Inst_RegFile_32x4__1342_/Q Inst_RegFile_32x4/_0459_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0466_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3/X ConfigBits\[344\]
+ ConfigBits\[345\] VGND VGND VPWR VPWR JS2BEG\[6\] sky130_fd_sc_hd__mux4_2
XFILLER_0_67_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1 net6 net24
+ net158 net211 ConfigBits\[286\] ConfigBits\[287\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XS4END_inbuf_4__0_ net187 VGND VGND VPWR VPWR S4BEG_i\[4\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput504 net504 VGND VGND VPWR VPWR WW4BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame5_bit1 net60 net96 VGND VGND VPWR VPWR ConfigBits\[223\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XW6END_inbuf_8__0_ net227 VGND VGND VPWR VPWR W6BEG_i\[8\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG2 net117 net17 net169
+ JS2BEG\[4\] ConfigBits\[170\] ConfigBits\[171\] VGND VGND VPWR VPWR J2MID_CDa_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XEE4BEG_outbuf_5__0_ EE4BEG_i\[5\] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 E2END[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1421_ net205 Inst_RegFile_32x4/_0073_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1421_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput345 net345 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput334 net334 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput378 net378 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput389 net389 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput367 net367 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput356 net356 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput323 net323 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1283_ Inst_RegFile_32x4/_0630_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0102_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput312 net312 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput301 net301 VGND VGND VPWR VPWR EE4BEG[9] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1352_ net205 Inst_RegFile_32x4/_0012_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1352_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0998_ Inst_RegFile_32x4__1391_/D Inst_RegFile_32x4__1391_/Q ConfigBits\[1\]
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0449_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG3 net114 net14 net166
+ net219 ConfigBits\[212\] ConfigBits\[213\] VGND VGND VPWR VPWR J2MID_EFb_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst0 net104
+ net156 net209 AD2 ConfigBits\[97\] ConfigBits\[98\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame12_bit22 net63 net84 VGND VGND VPWR VPWR ConfigBits\[20\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit11 net51 net84 VGND VGND VPWR VPWR ConfigBits\[9\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1 net24
+ net160 net182 net213 ConfigBits\[358\] ConfigBits\[359\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_13 J_l_GH_BEG\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0783_ Inst_RegFile_32x4__1426_/Q Inst_RegFile_32x4__1422_/Q Inst_RegFile_32x4/_0165_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0247_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0921_ Inst_RegFile_32x4/_0370_ Inst_RegFile_32x4/_0372_ Inst_RegFile_32x4/_0374_
+ Inst_RegFile_32x4/_0376_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0377_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_32x4__0852_ Inst_RegFile_32x4/_0309_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0310_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame2_bit4 net75 net93 VGND VGND VPWR VPWR ConfigBits\[322\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_46 JW2BEG\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_57 net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__1404_ net205 Inst_RegFile_32x4/_0056_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1404_/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_35 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 SS4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1266_ Inst_RegFile_32x4/_0620_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0095_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1335_ Inst_RegFile_32x4/_0659_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0125_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1197_ Inst_RegFile_32x4/_0577_ Inst_RegFile_32x4__1416_/Q Inst_RegFile_32x4/_0578_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput66 FrameData[25] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_8
Xinput55 FrameData[15] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0 net102
+ net110 net146 net2 ConfigBits\[270\] ConfigBits\[271\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
Xinput77 FrameData[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_8
Xinput22 E6END[10] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput44 EE4END[5] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput33 EE4END[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xinput11 E2END[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
XFILLER_0_24_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput88 FrameStrobe[16] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1120_ Inst_RegFile_32x4/_0473_ Inst_RegFile_32x4/_0513_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0534_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput99 FrameStrobe[8] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_16
XInst_RegFile_32x4__1051_ Inst_RegFile_32x4__1351_/Q Inst_RegFile_32x4/_0481_ Inst_RegFile_32x4/_0486_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0766_ Inst_RegFile_32x4/_0145_ Inst_RegFile_32x4/_0229_ Inst_RegFile_32x4/_0179_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0835_ Inst_RegFile_32x4__1356_/Q Inst_RegFile_32x4__1444_/Q Inst_RegFile_32x4/_0292_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0293_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0904_ Inst_RegFile_32x4__1369_/Q Inst_RegFile_32x4__1365_/Q Inst_RegFile_32x4/_0307_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0360_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame11_bit21 net62 net83 VGND VGND VPWR VPWR ConfigBits\[51\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame11_bit10 net50 net83 VGND VGND VPWR VPWR ConfigBits\[40\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0697_ Inst_RegFile_32x4/_0148_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0163_
+ sky130_fd_sc_hd__clkbuf_2
XSS4END_inbuf_11__0_ net195 VGND VGND VPWR VPWR SS4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1249_ Inst_RegFile_32x4/_0458_ Inst_RegFile_32x4/_0600_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0611_ sky130_fd_sc_hd__nand2_2
XInst_RegFile_32x4__1318_ Inst_RegFile_32x4/_0479_ Inst_RegFile_32x4__1466_/Q Inst_RegFile_32x4/_0647_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_outbuf_4__0_ FrameData_O_i\[4\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1 net159
+ net181 net212 net245 ConfigBits\[322\] ConfigBits\[323\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_inbuf_28__0_ net69 VGND VGND VPWR VPWR FrameData_O_i\[28\] sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1103_ Inst_RegFile_32x4/_0522_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0030_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1034_ Inst_RegFile_32x4/_0478_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0005_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0749_ Inst_RegFile_32x4/_0135_ Inst_RegFile_32x4/_0213_ Inst_RegFile_32x4/_0179_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0214_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0818_ Inst_RegFile_32x4/_0168_ Inst_RegFile_32x4/_0280_ Inst_RegFile_32x4/_0171_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0281_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XWW4END_inbuf_0__0_ net248 VGND VGND VPWR VPWR WW4BEG_i\[0\] sky130_fd_sc_hd__clkbuf_2
Xinput201 SS4END[6] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_19__0_ net59 VGND VGND VPWR VPWR FrameData_O_i\[19\] sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_7__0_ net98 VGND VGND VPWR VPWR FrameStrobe_O_i\[7\] sky130_fd_sc_hd__clkbuf_1
Xinput234 W6END[6] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_1
Xinput223 W2MID[5] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_2
Xinput212 W2END[2] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_4
Xinput245 WW4END[1] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_N4BEG3 net106 net121 net226 BD3 ConfigBits\[16\]
+ ConfigBits\[17\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__mux4_2
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame10_bit20 net61 net82 VGND VGND VPWR VPWR ConfigBits\[82\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit31 net73 net82 VGND VGND VPWR VPWR ConfigBits\[93\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst0 net102
+ net2 net154 AD0 ConfigBits\[47\] ConfigBits\[48\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1017_ Inst_RegFile_32x4/_0464_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0465_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2 net229
+ AD1 AD2 AD3 ConfigBits\[286\] ConfigBits\[287\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput505 net505 VGND VGND VPWR VPWR WW4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame5_bit2 net71 net96 VGND VGND VPWR VPWR ConfigBits\[224\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG3 net113 net165 net218
+ JW2BEG\[4\] ConfigBits\[172\] ConfigBits\[173\] VGND VGND VPWR VPWR J2MID_CDa_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XE6END_inbuf_0__0_ net25 VGND VGND VPWR VPWR E6BEG_i\[0\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_23_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 E2END[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1420_ net205 Inst_RegFile_32x4/_0072_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1420_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1351_ net205 Inst_RegFile_32x4/_0011_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1351_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput335 net335 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput346 net346 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput368 net368 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput357 net357 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput379 net379 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1282_ Inst_RegFile_32x4__1450_/Q Inst_RegFile_32x4/_0596_ Inst_RegFile_32x4/_0627_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0630_ sky130_fd_sc_hd__mux2_1
Xoutput313 net313 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput324 net324 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput302 net302 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0997_ Inst_RegFile_32x4/_0448_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1391_/D
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4END_inbuf_2__0_ net201 VGND VGND VPWR VPWR SS4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XEE4END_inbuf_11__0_ net39 VGND VGND VPWR VPWR EE4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst1 BD2 J2MID_ABa_BEG\[2\]
+ J2MID_CDa_BEG\[2\] J2END_EF_BEG\[2\] ConfigBits\[97\] ConfigBits\[98\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame12_bit23 net64 net84 VGND VGND VPWR VPWR ConfigBits\[21\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit12 net52 net84 VGND VGND VPWR VPWR ConfigBits\[10\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0920_ Inst_RegFile_32x4/_0296_ Inst_RegFile_32x4/_0375_ Inst_RegFile_32x4/_0340_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0376_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2 net229
+ AD0 AD1 AD3 ConfigBits\[358\] ConfigBits\[359\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
Xstrobe_outbuf_4__0_ FrameStrobe_O_i\[4\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_1
XANTENNA_14 N4BEG_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0782_ Inst_RegFile_32x4/_0239_ Inst_RegFile_32x4/_0241_ Inst_RegFile_32x4/_0243_
+ Inst_RegFile_32x4/_0245_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0246_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_32x4__0851_ B_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0309_ sky130_fd_sc_hd__inv_2
XANTENNA_25 SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_47 J_l_AB_BEG\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_ConfigMem_Inst_frame2_bit5 net76 net93 VGND VGND VPWR VPWR ConfigBits\[323\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_36 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__1334_ Inst_RegFile_32x4__1473_/Q Inst_RegFile_32x4/_0461_ Inst_RegFile_32x4/_0657_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_58 net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1403_ net205 Inst_RegFile_32x4/_0055_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1403_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1265_ Inst_RegFile_32x4__1443_/Q Inst_RegFile_32x4/_0598_ Inst_RegFile_32x4/_0616_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0620_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1196_ Inst_RegFile_32x4/_0554_ Inst_RegFile_32x4/_0571_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0578_ sky130_fd_sc_hd__nand2_2
XFILLER_0_69_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__1_/A1 ConfigBits\[82\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XEE4END_inbuf_1__0_ net44 VGND VGND VPWR VPWR EE4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_19__0_ net91 VGND VGND VPWR VPWR FrameStrobe_O_i\[19\] sky130_fd_sc_hd__clkbuf_2
XWW4BEG_outbuf_2__0_ WW4BEG_i\[2\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput67 FrameData[26] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_8
Xinput56 FrameData[16] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_8
Xinput78 FrameData[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1 net10
+ net154 net162 net207 ConfigBits\[270\] ConfigBits\[271\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xinput23 E6END[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 EE4END[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 EE4END[6] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput12 E2END[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XFILLER_0_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput89 FrameStrobe[17] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1050_ Inst_RegFile_32x4/_0489_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0010_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0903_ Inst_RegFile_32x4/_0334_ Inst_RegFile_32x4/_0358_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0359_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0765_ Inst_RegFile_32x4__1370_/Q Inst_RegFile_32x4__1366_/Q Inst_RegFile_32x4/_0177_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame11_bit11 net51 net83 VGND VGND VPWR VPWR ConfigBits\[41\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0834_ Inst_RegFile_32x4/_0291_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0292_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0696_ Inst_RegFile_32x4__1344_/Q Inst_RegFile_32x4__1392_/Q Inst_RegFile_32x4__1464_/Q
+ Inst_RegFile_32x4__1460_/Q Inst_RegFile_32x4/_0160_ Inst_RegFile_32x4/_0161_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0162_ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame11_bit22 net63 net83 VGND VGND VPWR VPWR ConfigBits\[52\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1317_ Inst_RegFile_32x4/_0649_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0117_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1248_ Inst_RegFile_32x4/_0610_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0087_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1179_ Inst_RegFile_32x4/_0567_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0061_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XE6BEG_outbuf_5__0_ E6BEG_i\[5\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0 net104
+ net112 net4 net12 ConfigBits\[310\] ConfigBits\[311\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2 net226
+ AD0 AD2 AD3 ConfigBits\[322\] ConfigBits\[323\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XN4END_inbuf_4__0_ net135 VGND VGND VPWR VPWR N4BEG_i\[4\] sky130_fd_sc_hd__buf_2
XFILLER_0_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1102_ Inst_RegFile_32x4__1370_/Q Inst_RegFile_32x4/_0498_ Inst_RegFile_32x4/_0519_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0522_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1033_ Inst_RegFile_32x4__1345_/Q Inst_RegFile_32x4/_0477_ Inst_RegFile_32x4/_0475_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0478_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame8_bit0 net49 net99 VGND VGND VPWR VPWR ConfigBits\[126\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0748_ Inst_RegFile_32x4__1433_/Q Inst_RegFile_32x4__1429_/Q Inst_RegFile_32x4/_0177_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0213_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0817_ Inst_RegFile_32x4__1419_/Q Inst_RegFile_32x4__1415_/Q Inst_RegFile_32x4/_0169_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0280_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0679_ Inst_RegFile_32x4/_0134_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0145_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput202 SS4END[7] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
Xinput235 W6END[7] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
Xinput224 W2MID[6] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_4
Xinput213 W2END[3] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_4
Xinput246 WW4END[2] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame10_bit21 net62 net82 VGND VGND VPWR VPWR ConfigBits\[83\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit10 net50 net82 VGND VGND VPWR VPWR ConfigBits\[72\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst1 BD0 J2MID_EFa_BEG\[2\]
+ J2MID_GHa_BEG\[2\] J2END_AB_BEG\[0\] ConfigBits\[47\] ConfigBits\[48\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_cus_mux41_buf_inst0 net107 net159
+ J2MID_ABa_BEG\[1\] J2MID_ABb_BEG\[2\] ConfigBits\[133\] ConfigBits\[134\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1016_ D2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0464_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[286\] ConfigBits\[287\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput506 net506 VGND VGND VPWR VPWR WW4BEG[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame5_bit3 net74 net96 VGND VGND VPWR VPWR ConfigBits\[225\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput325 net325 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__clkbuf_4
Xoutput314 net314 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput303 net303 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1350_ net205 Inst_RegFile_32x4/_0010_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1350_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput336 net336 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput347 net347 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XNN4BEG_outbuf_5__0_ NN4BEG_i\[5\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_1
Xoutput369 net369 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput358 net358 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1281_ Inst_RegFile_32x4/_0629_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0101_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XN4BEG_outbuf_9__0_ N4BEG_i\[9\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0996_ Inst_RegFile_32x4/_0426_ Inst_RegFile_32x4/_0432_ Inst_RegFile_32x4/_0441_
+ Inst_RegFile_32x4/_0447_ B_ADR3 B_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0448_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSS4BEG_outbuf_8__0_ SS4BEG_i\[8\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame12_bit24 net65 net84 VGND VGND VPWR VPWR ConfigBits\[22\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit13 net53 net84 VGND VGND VPWR VPWR ConfigBits\[11\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix__49_ JW2BEG\[1\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[358\] ConfigBits\[359\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_15 N4BEG_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0781_ Inst_RegFile_32x4/_0135_ Inst_RegFile_32x4/_0244_ Inst_RegFile_32x4/_0179_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0245_ sky130_fd_sc_hd__a21o_1
XANTENNA_37 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0850_ Inst_RegFile_32x4__1368_/Q Inst_RegFile_32x4__1364_/Q Inst_RegFile_32x4/_0307_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0308_ sky130_fd_sc_hd__mux2_1
XANTENNA_26 SS4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_ConfigMem_Inst_frame2_bit6 net77 net93 VGND VGND VPWR VPWR ConfigBits\[324\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_48 J_l_AB_BEG\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1264_ Inst_RegFile_32x4/_0619_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0094_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1333_ Inst_RegFile_32x4/_0658_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0124_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0 net101
+ net105 net1 net5 ConfigBits\[346\] ConfigBits\[347\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1402_ net205 Inst_RegFile_32x4/_0054_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1402_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1195_ Inst_RegFile_32x4/_0450_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0577_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_ConfigMem_Inst_frame12_bit2 net71 net84 VGND VGND VPWR VPWR ConfigBits\[0\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XW6BEG_outbuf_9__0_ W6BEG_i\[9\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0979_ Inst_RegFile_32x4__1347_/Q Inst_RegFile_32x4__1395_/Q Inst_RegFile_32x4__1467_/Q
+ Inst_RegFile_32x4__1463_/Q Inst_RegFile_32x4/_0307_ Inst_RegFile_32x4/_0295_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0431_ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2 net209
+ AD0 AD1 AD2 ConfigBits\[270\] ConfigBits\[271\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput13 E2MID[0] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput68 FrameData[27] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_6
Xinput57 FrameData[17] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_8
Xinput79 FrameData[8] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_4
Xinput24 E6END[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_4
Xinput35 EE4END[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
Xinput46 EE4END[7] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XNN4END_inbuf_2__0_ net149 VGND VGND VPWR VPWR NN4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0833_ B_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0291_ sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__0902_ Inst_RegFile_32x4__1377_/Q Inst_RegFile_32x4__1373_/Q Inst_RegFile_32x4/_0303_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0358_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame11_bit23 net64 net83 VGND VGND VPWR VPWR ConfigBits\[53\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame11_bit12 net52 net83 VGND VGND VPWR VPWR ConfigBits\[42\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0764_ Inst_RegFile_32x4/_0173_ Inst_RegFile_32x4/_0227_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0228_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0695_ A_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0161_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1247_ Inst_RegFile_32x4/_0584_ Inst_RegFile_32x4__1435_/Q Inst_RegFile_32x4/_0606_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0610_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1316_ Inst_RegFile_32x4/_0477_ Inst_RegFile_32x4__1465_/Q Inst_RegFile_32x4/_0647_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1178_ Inst_RegFile_32x4/_0462_ Inst_RegFile_32x4__1409_/Q Inst_RegFile_32x4/_0565_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_29__0_ FrameData_O_i\[29\] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1 net40
+ net154 net156 net164 ConfigBits\[310\] ConfigBits\[311\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[322\] ConfigBits\[323\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1101_ Inst_RegFile_32x4/_0521_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0029_
+ sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_9__0_ S4BEG_i\[9\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame8_bit1 net60 net99 VGND VGND VPWR VPWR ConfigBits\[127\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1032_ D1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0477_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0816_ Inst_RegFile_32x4/_0182_ Inst_RegFile_32x4/_0278_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0279_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0747_ Inst_RegFile_32x4/_0173_ Inst_RegFile_32x4/_0211_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0212_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0678_ Inst_RegFile_32x4/_0141_ Inst_RegFile_32x4/_0143_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0144_ sky130_fd_sc_hd__and2b_1
Xinput203 SS4END[8] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
Xinput236 W6END[8] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_1
Xinput247 WW4END[3] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__buf_2
Xinput225 W2MID[7] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_2
Xinput214 W2END[4] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XS4END_inbuf_7__0_ net175 VGND VGND VPWR VPWR S4BEG_i\[7\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame10_bit22 net63 net82 VGND VGND VPWR VPWR ConfigBits\[84\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit11 net51 net82 VGND VGND VPWR VPWR ConfigBits\[73\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_cus_mux41_buf_inst1 J2END_EF_BEG\[3\]
+ JN2BEG\[6\] JS2BEG\[6\] JW2BEG\[6\] ConfigBits\[133\] ConfigBits\[134\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1015_ Inst_RegFile_32x4/_0463_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0001_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XEE4BEG_outbuf_8__0_ EE4BEG_i\[8\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3/X ConfigBits\[288\]
+ ConfigBits\[289\] VGND VGND VPWR VPWR JE2BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_W1BEG0 BD1 J2MID_CDb_BEG\[3\] JS2BEG\[3\]
+ J_l_CD_BEG\[1\] ConfigBits\[86\] ConfigBits\[87\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__mux4_1
XFILLER_0_66_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame5_bit4 net75 net96 VGND VGND VPWR VPWR ConfigBits\[226\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput359 net359 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput348 net348 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput337 net337 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput326 net326 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1280_ Inst_RegFile_32x4__1449_/Q Inst_RegFile_32x4/_0594_ Inst_RegFile_32x4/_0627_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0629_ sky130_fd_sc_hd__mux2_1
Xoutput315 net315 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__clkbuf_4
Xoutput304 net304 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0995_ Inst_RegFile_32x4/_0443_ Inst_RegFile_32x4/_0445_ Inst_RegFile_32x4/_0446_
+ Inst_RegFile_32x4/_0324_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0447_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame12_bit25 net66 net84 VGND VGND VPWR VPWR ConfigBits\[23\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit14 net54 net84 VGND VGND VPWR VPWR ConfigBits\[12\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix__48_ JW2BEG\[0\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3/X ConfigBits\[360\]
+ ConfigBits\[361\] VGND VGND VPWR VPWR JW2BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_16 N4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__0780_ Inst_RegFile_32x4__1434_/Q Inst_RegFile_32x4__1430_/Q Inst_RegFile_32x4/_0177_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0244_ sky130_fd_sc_hd__mux2_1
XANTENNA_27 W6BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_ConfigMem_Inst_frame2_bit7 net78 net93 VGND VGND VPWR VPWR ConfigBits\[325\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_49 J_l_AB_BEG\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__1401_ net205 Inst_RegFile_32x4/_0053_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1401_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1263_ Inst_RegFile_32x4__1442_/Q Inst_RegFile_32x4/_0596_ Inst_RegFile_32x4/_0616_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0619_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1332_ Inst_RegFile_32x4__1472_/Q Inst_RegFile_32x4/_0450_ Inst_RegFile_32x4/_0657_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0658_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1 net153
+ net157 net189 net206 ConfigBits\[346\] ConfigBits\[347\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1194_ Inst_RegFile_32x4/_0576_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0067_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame12_bit3 net74 net84 VGND VGND VPWR VPWR ConfigBits\[1\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XNN4END_inbuf_11__0_ net143 VGND VGND VPWR VPWR NN4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0978_ Inst_RegFile_32x4/_0302_ Inst_RegFile_32x4/_0429_ B_ADR2
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0430_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_12__0_ FrameStrobe_O_i\[12\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3 AD3 BD1
+ BD2 BD3 ConfigBits\[270\] ConfigBits\[271\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput25 E6END[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 EE4END[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput14 E2MID[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput69 FrameData[28] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_6
Xinput58 FrameData[18] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_8
Xdata_outbuf_7__0_ FrameData_O_i\[7\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_1
Xinput47 EE4END[8] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0763_ Inst_RegFile_32x4__1378_/Q Inst_RegFile_32x4__1374_/Q Inst_RegFile_32x4/_0142_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0227_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0901_ Inst_RegFile_32x4/_0296_ Inst_RegFile_32x4/_0356_ Inst_RegFile_32x4/_0300_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0357_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0832_ Inst_RegFile_32x4/_0289_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0290_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_70_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame11_bit24 net65 net83 VGND VGND VPWR VPWR ConfigBits\[54\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame11_bit13 net53 net83 VGND VGND VPWR VPWR ConfigBits\[43\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0694_ Inst_RegFile_32x4/_0136_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0160_
+ sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1246_ Inst_RegFile_32x4/_0609_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0086_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1315_ Inst_RegFile_32x4/_0648_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0116_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1177_ Inst_RegFile_32x4/_0566_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0060_
+ sky130_fd_sc_hd__clkbuf_1
XWW4END_inbuf_3__0_ net251 VGND VGND VPWR VPWR WW4BEG_i\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2 net209
+ AD0 AD1 AD2 ConfigBits\[310\] ConfigBits\[311\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3/X ConfigBits\[324\]
+ ConfigBits\[325\] VGND VGND VPWR VPWR JS2BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1100_ Inst_RegFile_32x4__1369_/Q Inst_RegFile_32x4/_0496_ Inst_RegFile_32x4/_0519_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0521_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1031_ Inst_RegFile_32x4/_0476_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0004_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame8_bit2 net71 net99 VGND VGND VPWR VPWR ConfigBits\[128\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0746_ Inst_RegFile_32x4__1441_/Q Inst_RegFile_32x4__1437_/Q Inst_RegFile_32x4/_0174_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0211_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0815_ Inst_RegFile_32x4__1427_/Q Inst_RegFile_32x4__1423_/Q Inst_RegFile_32x4/_0165_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0677_ Inst_RegFile_32x4__1376_/Q Inst_RegFile_32x4__1372_/Q Inst_RegFile_32x4/_0142_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0143_ sky130_fd_sc_hd__mux2_1
Xinput204 SS4END[9] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1229_ Inst_RegFile_32x4/_0599_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0079_
+ sky130_fd_sc_hd__clkbuf_1
Xinput226 W6END[0] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_4
Xinput237 W6END[9] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_1
Xinput248 WW4END[4] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput215 W2END[5] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame10_bit23 net64 net82 VGND VGND VPWR VPWR ConfigBits\[85\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit12 net52 net82 VGND VGND VPWR VPWR ConfigBits\[74\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1014_ Inst_RegFile_32x4/_0462_ Inst_RegFile_32x4__1341_/Q Inst_RegFile_32x4/_0459_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0729_ Inst_RegFile_32x4__1405_/Q Inst_RegFile_32x4__1381_/Q Inst_RegFile_32x4/_0137_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XE6END_inbuf_3__0_ net28 VGND VGND VPWR VPWR E6BEG_i\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_W1BEG1 BD2 J2MID_EFb_BEG\[0\] JS2BEG\[0\]
+ J_l_EF_BEG\[2\] ConfigBits\[88\] ConfigBits\[89\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__mux4_1
XFILLER_0_66_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame9_bit30 net72 net100 VGND VGND VPWR VPWR ConfigBits\[124\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame5_bit5 net76 net96 VGND VGND VPWR VPWR ConfigBits\[227\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4END_inbuf_5__0_ net204 VGND VGND VPWR VPWR SS4BEG_i\[5\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput349 net349 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput338 net338 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput316 net316 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__clkbuf_4
Xoutput305 net305 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput327 net327 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_7__0_ FrameStrobe_O_i\[7\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0994_ Inst_RegFile_32x4__1411_/Q Inst_RegFile_32x4__1343_/Q Inst_RegFile_32x4__1403_/Q
+ Inst_RegFile_32x4__1471_/Q Inst_RegFile_32x4/_0321_ Inst_RegFile_32x4/_0322_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0446_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame12_bit26 net67 net84 VGND VGND VPWR VPWR ConfigBits\[24\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit15 net55 net84 VGND VGND VPWR VPWR ConfigBits\[13\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__47_ net172 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkbuf_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XEE4END_inbuf_4__0_ net47 VGND VGND VPWR VPWR EE4BEG_i\[4\] sky130_fd_sc_hd__clkbuf_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_inbuf_1__0_ net60 VGND VGND VPWR VPWR FrameData_O_i\[1\] sky130_fd_sc_hd__buf_1
XFILLER_0_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame2_bit8 net79 net93 VGND VGND VPWR VPWR ConfigBits\[326\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XWW4BEG_outbuf_5__0_ WW4BEG_i\[5\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_1
XANTENNA_17 NN4BEG_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_39 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_32x4__1400_ net205 Inst_RegFile_32x4/_0052_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1400_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1262_ Inst_RegFile_32x4/_0618_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0093_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1193_ Inst_RegFile_32x4/_0468_ Inst_RegFile_32x4__1415_/Q Inst_RegFile_32x4/_0572_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0576_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2 net208
+ AD0 AD1 AD2 ConfigBits\[346\] ConfigBits\[347\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1331_ Inst_RegFile_32x4/_0485_ Inst_RegFile_32x4/_0626_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0657_ sky130_fd_sc_hd__nor2_2
XFILLER_0_2_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame12_bit4 net75 net84 VGND VGND VPWR VPWR ConfigBits\[2\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0977_ Inst_RegFile_32x4__1355_/Q Inst_RegFile_32x4__1351_/Q Inst_RegFile_32x4/_0303_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput59 FrameData[19] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3/X ConfigBits\[272\]
+ ConfigBits\[273\] VGND VGND VPWR VPWR JN2BEG\[4\] sky130_fd_sc_hd__mux4_2
Xinput26 E6END[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 EE4END[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput48 EE4END[9] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
Xinput15 E2MID[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XE6BEG_outbuf_8__0_ E6BEG_i\[8\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0900_ Inst_RegFile_32x4__1405_/Q Inst_RegFile_32x4__1381_/Q Inst_RegFile_32x4/_0298_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0762_ Inst_RegFile_32x4/_0185_ Inst_RegFile_32x4/_0225_ Inst_RegFile_32x4/_0139_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0226_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0831_ B_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0289_ sky130_fd_sc_hd__buf_1
XFILLER_0_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame11_bit25 net66 net83 VGND VGND VPWR VPWR ConfigBits\[55\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame11_bit14 net54 net83 VGND VGND VPWR VPWR ConfigBits\[44\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0693_ Inst_RegFile_32x4/_0141_ Inst_RegFile_32x4/_0157_ Inst_RegFile_32x4/_0158_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0159_ sky130_fd_sc_hd__a21o_1
XN4END_inbuf_7__0_ net123 VGND VGND VPWR VPWR N4BEG_i\[7\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1314_ Inst_RegFile_32x4/_0470_ Inst_RegFile_32x4__1464_/Q Inst_RegFile_32x4/_0647_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1245_ Inst_RegFile_32x4/_0582_ Inst_RegFile_32x4__1434_/Q Inst_RegFile_32x4/_0606_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0609_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1176_ Inst_RegFile_32x4/_0451_ Inst_RegFile_32x4__1408_/Q Inst_RegFile_32x4/_0565_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3 AD3 BD0
+ BD1 BD3 ConfigBits\[310\] ConfigBits\[311\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1030_ Inst_RegFile_32x4__1344_/Q Inst_RegFile_32x4/_0470_ Inst_RegFile_32x4/_0475_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame8_bit3 net74 net99 VGND VGND VPWR VPWR ConfigBits\[129\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0814_ Inst_RegFile_32x4/_0270_ Inst_RegFile_32x4/_0272_ Inst_RegFile_32x4/_0274_
+ Inst_RegFile_32x4/_0276_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0277_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_32x4__0745_ Inst_RegFile_32x4/_0168_ Inst_RegFile_32x4/_0209_ Inst_RegFile_32x4/_0171_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0210_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0676_ Inst_RegFile_32x4/_0130_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0142_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1228_ Inst_RegFile_32x4__1427_/Q Inst_RegFile_32x4/_0598_ Inst_RegFile_32x4/_0592_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0599_ sky130_fd_sc_hd__mux2_1
Xinput227 W6END[10] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1159_ Inst_RegFile_32x4/_0556_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0052_
+ sky130_fd_sc_hd__clkbuf_1
Xinput249 WW4END[5] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_1
Xinput205 UserCLK VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_16
Xinput216 W2END[6] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
Xinput238 WW4END[0] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_2
XFILLER_0_19_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame10_bit13 net53 net82 VGND VGND VPWR VPWR ConfigBits\[75\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit24 net65 net82 VGND VGND VPWR VPWR ConfigBits\[86\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1013_ Inst_RegFile_32x4/_0461_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0462_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0728_ Inst_RegFile_32x4/_0129_ Inst_RegFile_32x4/_0192_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0193_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_W1BEG2 BD3 J2MID_GHb_BEG\[1\] JS2BEG\[1\]
+ J_l_GH_BEG\[3\] ConfigBits\[90\] ConfigBits\[91\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame9_bit31 net73 net100 VGND VGND VPWR VPWR ConfigBits\[125\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit20 net61 net100 VGND VGND VPWR VPWR ConfigBits\[114\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame5_bit6 net77 net96 VGND VGND VPWR VPWR ConfigBits\[228\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XNN4BEG_outbuf_8__0_ NN4BEG_i\[8\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__63_ net225 VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_10__0_ FrameData_O_i\[10\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput339 net339 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput317 net317 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__clkbuf_4
Xoutput306 net306 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput328 net328 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0993_ Inst_RegFile_32x4/_0329_ Inst_RegFile_32x4/_0444_ Inst_RegFile_32x4/_0332_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__46_ net171 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame12_bit27 net68 net84 VGND VGND VPWR VPWR ConfigBits\[25\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit16 net56 net84 VGND VGND VPWR VPWR ConfigBits\[14\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit30 net72 net99 VGND VGND VPWR VPWR ConfigBits\[156\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_18 NN4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RegFile_ConfigMem_Inst_frame2_bit9 net80 net93 VGND VGND VPWR VPWR ConfigBits\[327\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1330_ Inst_RegFile_32x4/_0656_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0123_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1261_ Inst_RegFile_32x4__1441_/Q Inst_RegFile_32x4/_0594_ Inst_RegFile_32x4/_0616_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1192_ Inst_RegFile_32x4/_0575_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0066_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3 AD3 BD0
+ BD1 BD2 ConfigBits\[346\] ConfigBits\[347\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XW6END_inbuf_1__0_ net231 VGND VGND VPWR VPWR W6BEG_i\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XNN4END_inbuf_5__0_ net152 VGND VGND VPWR VPWR NN4BEG_i\[5\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0 net101
+ net107 net129 net144 ConfigBits\[290\] ConfigBits\[291\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame12_bit5 net76 net84 VGND VGND VPWR VPWR ConfigBits\[3\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0976_ Inst_RegFile_32x4/_0349_ Inst_RegFile_32x4/_0427_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0428_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__1459_ net205 Inst_RegFile_32x4/_0111_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1459_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix__29_ net118 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_1
XFILLER_0_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 FrameData[0] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_4
Xinput27 E6END[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput38 EE4END[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput16 E2MID[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XWW4END_inbuf_11__0_ net244 VGND VGND VPWR VPWR WW4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0830_ Inst_RegFile_32x4/_0288_ VGND VGND VPWR VPWR AD3 sky130_fd_sc_hd__buf_12
XInst_RegFile_32x4__0761_ Inst_RegFile_32x4__1406_/Q Inst_RegFile_32x4__1382_/Q Inst_RegFile_32x4/_0137_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0692_ A_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0158_ sky130_fd_sc_hd__buf_2
XInst_RegFile_ConfigMem_Inst_frame11_bit26 net67 net83 VGND VGND VPWR VPWR ConfigBits\[56\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame11_bit15 net55 net83 VGND VGND VPWR VPWR ConfigBits\[45\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1244_ Inst_RegFile_32x4/_0608_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0085_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1313_ Inst_RegFile_32x4/_0471_ Inst_RegFile_32x4/_0554_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0647_ sky130_fd_sc_hd__nand2_2
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1175_ Inst_RegFile_32x4/_0455_ Inst_RegFile_32x4/_0474_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0565_ sky130_fd_sc_hd__nand2_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG0 net146 net11 net163 net216
+ ConfigBits\[230\] ConfigBits\[231\] VGND VGND VPWR VPWR J2END_CD_BEG\[0\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0959_ Inst_RegFile_32x4/_0346_ Inst_RegFile_32x4/_0412_ Inst_RegFile_32x4/_0332_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0413_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3/X ConfigBits\[312\]
+ ConfigBits\[313\] VGND VGND VPWR VPWR JE2BEG\[6\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst0 net103
+ net3 net208 AD1 ConfigBits\[18\] ConfigBits\[19\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0813_ Inst_RegFile_32x4/_0135_ Inst_RegFile_32x4/_0275_ Inst_RegFile_32x4/_0148_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame8_bit4 net75 net99 VGND VGND VPWR VPWR ConfigBits\[130\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0744_ Inst_RegFile_32x4__1449_/Q Inst_RegFile_32x4__1473_/Q Inst_RegFile_32x4/_0156_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0675_ Inst_RegFile_32x4/_0128_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0141_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1227_ D3 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0598_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput206 W1END[0] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_4
Xinput217 W2END[7] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput228 W6END[11] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1089_ Inst_RegFile_32x4__1364_/Q Inst_RegFile_32x4/_0491_ Inst_RegFile_32x4/_0514_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0515_ sky130_fd_sc_hd__mux2_1
Xinput239 WW4END[10] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1158_ Inst_RegFile_32x4/_0451_ Inst_RegFile_32x4__1400_/Q Inst_RegFile_32x4/_0555_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0 net103
+ net109 net146 net9 ConfigBits\[362\] ConfigBits\[363\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame10_bit25 net66 net82 VGND VGND VPWR VPWR ConfigBits\[87\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit14 net54 net82 VGND VGND VPWR VPWR ConfigBits\[76\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1012_ D1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0461_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0727_ Inst_RegFile_32x4__1357_/Q Inst_RegFile_32x4__1445_/Q Inst_RegFile_32x4/_0131_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_inbuf_30__0_ net72 VGND VGND VPWR VPWR FrameData_O_i\[30\] sky130_fd_sc_hd__buf_1
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame9_bit21 net62 net100 VGND VGND VPWR VPWR ConfigBits\[115\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit10 net50 net100 VGND VGND VPWR VPWR ConfigBits\[104\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_W1BEG3 AD0 J2MID_ABb_BEG\[2\] JS2BEG\[2\]
+ J_l_AB_BEG\[0\] ConfigBits\[92\] ConfigBits\[93\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__mux4_1
Xdata_inbuf_21__0_ net62 VGND VGND VPWR VPWR FrameData_O_i\[21\] sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__1_/A1 ConfigBits\[40\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame5_bit7 net78 net96 VGND VGND VPWR VPWR ConfigBits\[229\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix__62_ net224 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_0__0_ net81 VGND VGND VPWR VPWR FrameStrobe_O_i\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_inbuf_12__0_ net52 VGND VGND VPWR VPWR FrameData_O_i\[12\] sky130_fd_sc_hd__buf_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0 net144
+ net4 net196 net209 ConfigBits\[106\] ConfigBits\[107\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0 net108
+ net2 net8 net41 ConfigBits\[326\] ConfigBits\[327\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput307 net307 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput318 net318 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__clkbuf_4
Xoutput329 net329 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0992_ Inst_RegFile_32x4__1419_/Q Inst_RegFile_32x4__1415_/Q Inst_RegFile_32x4/_0330_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1475_ net205 Inst_RegFile_32x4/_0127_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1475_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame12_bit28 net69 net84 VGND VGND VPWR VPWR ConfigBits\[26\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit17 net57 net84 VGND VGND VPWR VPWR ConfigBits\[15\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__45_ net170 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit20 net61 net99 VGND VGND VPWR VPWR ConfigBits\[146\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame8_bit31 net73 net99 VGND VGND VPWR VPWR ConfigBits\[157\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_15__0_ FrameStrobe_O_i\[15\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_1
XANTENNA_19 NN4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1260_ Inst_RegFile_32x4/_0617_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0092_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3/X ConfigBits\[348\]
+ ConfigBits\[349\] VGND VGND VPWR VPWR JS2BEG\[7\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__1191_ Inst_RegFile_32x4/_0465_ Inst_RegFile_32x4__1414_/Q Inst_RegFile_32x4/_0572_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0575_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame12_bit6 net77 net84 VGND VGND VPWR VPWR ConfigBits\[4\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1 net7 net21
+ net159 net212 ConfigBits\[290\] ConfigBits\[291\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0975_ Inst_RegFile_32x4__1363_/Q Inst_RegFile_32x4__1399_/Q Inst_RegFile_32x4/_0297_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1458_ net205 Inst_RegFile_32x4/_0110_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1458_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1389_ net205 Inst_RegFile_32x4__1389_/D VGND VGND VPWR VPWR Inst_RegFile_32x4__1389_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__28_ net117 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_1
XWW4END_inbuf_6__0_ net239 VGND VGND VPWR VPWR WW4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_2
Xinput28 E6END[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 EE4END[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
Xinput17 E2MID[4] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame11_bit27 net68 net83 VGND VGND VPWR VPWR ConfigBits\[57\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame11_bit16 net56 net83 VGND VGND VPWR VPWR ConfigBits\[46\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0760_ Inst_RegFile_32x4/_0129_ Inst_RegFile_32x4/_0223_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0224_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0691_ Inst_RegFile_32x4__1352_/Q Inst_RegFile_32x4__1348_/Q Inst_RegFile_32x4/_0156_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0157_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1243_ Inst_RegFile_32x4/_0580_ Inst_RegFile_32x4__1433_/Q Inst_RegFile_32x4/_0606_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1312_ Inst_RegFile_32x4/_0646_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0115_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1174_ Inst_RegFile_32x4/_0564_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0059_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame7_bit30 net72 net98 VGND VGND VPWR VPWR ConfigBits\[188\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0958_ Inst_RegFile_32x4__1418_/Q Inst_RegFile_32x4__1414_/Q Inst_RegFile_32x4/_0330_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0412_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG1 net107 net7 net159 net246
+ ConfigBits\[232\] ConfigBits\[233\] VGND VGND VPWR VPWR J2END_CD_BEG\[1\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__0889_ Inst_RegFile_32x4__1416_/Q Inst_RegFile_32x4__1412_/Q Inst_RegFile_32x4/_0330_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0347_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__1_/A1 ConfigBits\[23\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
Xoutput490 net490 VGND VGND VPWR VPWR W6BEG[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst1 BD1 J2MID_ABb_BEG\[1\]
+ J2MID_CDb_BEG\[1\] J2END_GH_BEG\[1\] ConfigBits\[18\] ConfigBits\[19\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst0 net101
+ net153 net206 AD3 ConfigBits\[100\] ConfigBits\[101\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame8_bit5 net76 net99 VGND VGND VPWR VPWR ConfigBits\[131\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0812_ Inst_RegFile_32x4__1435_/Q Inst_RegFile_32x4__1431_/Q Inst_RegFile_32x4/_0137_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0743_ Inst_RegFile_32x4/_0152_ Inst_RegFile_32x4/_0207_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0208_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0674_ Inst_RegFile_32x4/_0135_ Inst_RegFile_32x4/_0138_ Inst_RegFile_32x4/_0139_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0140_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__1226_ Inst_RegFile_32x4/_0597_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0078_
+ sky130_fd_sc_hd__clkbuf_1
Xinput229 W6END[1] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_4
XInst_RegFile_32x4__1157_ Inst_RegFile_32x4/_0455_ Inst_RegFile_32x4/_0554_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0555_ sky130_fd_sc_hd__nand2_2
Xinput207 W1END[1] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_4
Xinput218 W2MID[0] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1088_ Inst_RegFile_32x4/_0485_ Inst_RegFile_32x4/_0513_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0514_ sky130_fd_sc_hd__nor2_2
XFILLER_0_66_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1 net21
+ net161 net173 net214 ConfigBits\[362\] ConfigBits\[363\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xstrobe_inbuf_12__0_ net84 VGND VGND VPWR VPWR FrameStrobe_O_i\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XE6END_inbuf_6__0_ net31 VGND VGND VPWR VPWR E6BEG_i\[6\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame10_bit26 net67 net82 VGND VGND VPWR VPWR ConfigBits\[88\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit15 net55 net82 VGND VGND VPWR VPWR ConfigBits\[77\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1011_ Inst_RegFile_32x4/_0460_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0000_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0726_ Inst_RegFile_32x4/_0191_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1384_/D
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0 net103
+ net111 net145 net3 ConfigBits\[274\] ConfigBits\[275\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1209_ Inst_RegFile_32x4/_0577_ Inst_RegFile_32x4__1420_/Q Inst_RegFile_32x4/_0586_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0587_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG0 net130 net33 net182 JN2BEG\[4\]
+ ConfigBits\[406\] ConfigBits\[407\] VGND VGND VPWR VPWR J_l_GH_BEG\[0\] sky130_fd_sc_hd__mux4_1
XSS4END_inbuf_8__0_ net192 VGND VGND VPWR VPWR SS4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame9_bit22 net63 net100 VGND VGND VPWR VPWR ConfigBits\[116\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit11 net51 net100 VGND VGND VPWR VPWR ConfigBits\[105\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame5_bit8 net79 net96 VGND VGND VPWR VPWR ConfigBits\[230\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst0 net103
+ net3 net208 AD1 ConfigBits\[74\] ConfigBits\[75\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix__61_ net223 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__0709_ Inst_RegFile_32x4__1440_/Q Inst_RegFile_32x4__1436_/Q Inst_RegFile_32x4/_0174_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1 AD0 AD1
+ AD2 AD3 ConfigBits\[106\] ConfigBits\[107\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1 net24
+ net160 net182 net213 ConfigBits\[326\] ConfigBits\[327\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XEE4END_inbuf_7__0_ net35 VGND VGND VPWR VPWR EE4BEG_i\[7\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput319 net319 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__clkbuf_4
Xoutput308 net308 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_inbuf_4__0_ net75 VGND VGND VPWR VPWR FrameData_O_i\[4\] sky130_fd_sc_hd__buf_1
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0991_ Inst_RegFile_32x4/_0343_ Inst_RegFile_32x4/_0442_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0443_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XWW4BEG_outbuf_8__0_ WW4BEG_i\[8\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1474_ net205 Inst_RegFile_32x4/_0126_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1474_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__1_/A1 ConfigBits\[102\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame12_bit29 net70 net84 VGND VGND VPWR VPWR ConfigBits\[27\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame12_bit18 net58 net84 VGND VGND VPWR VPWR ConfigBits\[16\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__44_ net169 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame8_bit10 net50 net99 VGND VGND VPWR VPWR ConfigBits\[136\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit21 net62 net99 VGND VGND VPWR VPWR ConfigBits\[147\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1190_ Inst_RegFile_32x4/_0574_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0065_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2 net226
+ AD0 AD2 AD3 ConfigBits\[290\] ConfigBits\[291\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame12_bit7 net78 net84 VGND VGND VPWR VPWR ConfigBits\[5\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0974_ Inst_RegFile_32x4/_0419_ Inst_RegFile_32x4/_0421_ Inst_RegFile_32x4/_0423_
+ Inst_RegFile_32x4/_0425_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0426_ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1457_ net205 Inst_RegFile_32x4/_0109_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1457_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1388_ net205 Inst_RegFile_32x4__1388_/D VGND VGND VPWR VPWR Inst_RegFile_32x4__1388_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix__27_ net116 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 E2MID[5] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame1_bit0 net49 net92 VGND VGND VPWR VPWR ConfigBits\[350\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput29 E6END[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG0 net120 net20 net172
+ net225 ConfigBits\[214\] ConfigBits\[215\] VGND VGND VPWR VPWR J2MID_GHb_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XN4BEG_outbuf_2__0_ N4BEG_i\[2\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame11_bit17 net57 net83 VGND VGND VPWR VPWR ConfigBits\[47\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0690_ Inst_RegFile_32x4/_0130_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0156_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame11_bit28 net69 net83 VGND VGND VPWR VPWR ConfigBits\[58\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1242_ Inst_RegFile_32x4/_0607_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0084_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1173_ Inst_RegFile_32x4__1407_/Q Inst_RegFile_32x4/_0532_ Inst_RegFile_32x4/_0560_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0564_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame7_bit20 net61 net98 VGND VGND VPWR VPWR ConfigBits\[178\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1311_ Inst_RegFile_32x4/_0481_ Inst_RegFile_32x4__1463_/Q Inst_RegFile_32x4/_0642_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0646_ sky130_fd_sc_hd__mux2_1
XSS4BEG_outbuf_1__0_ SS4BEG_i\[1\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame7_bit31 net73 net98 VGND VGND VPWR VPWR ConfigBits\[189\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0888_ Inst_RegFile_32x4/_0295_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0346_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_32x4__0957_ Inst_RegFile_32x4/_0343_ Inst_RegFile_32x4/_0410_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0411_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG2 net109 net9 net197 net214
+ ConfigBits\[234\] ConfigBits\[235\] VGND VGND VPWR VPWR J2END_CD_BEG\[2\] sky130_fd_sc_hd__mux4_2
Xoutput480 net480 VGND VGND VPWR VPWR W6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput491 net491 VGND VGND VPWR VPWR WW4BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst1 BD3 J2MID_EFb_BEG\[1\]
+ J2MID_GHb_BEG\[1\] J2END_CD_BEG\[2\] ConfigBits\[100\] ConfigBits\[101\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XW6BEG_outbuf_2__0_ W6BEG_i\[2\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame8_bit6 net77 net99 VGND VGND VPWR VPWR ConfigBits\[132\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0811_ Inst_RegFile_32x4/_0129_ Inst_RegFile_32x4/_0273_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0274_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0742_ Inst_RegFile_32x4__1457_/Q Inst_RegFile_32x4__1453_/Q Inst_RegFile_32x4/_0165_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0673_ A_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0139_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1225_ Inst_RegFile_32x4__1426_/Q Inst_RegFile_32x4/_0596_ Inst_RegFile_32x4/_0592_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0597_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1156_ Inst_RegFile_32x4/_0484_ Inst_RegFile_32x4/_0492_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0554_ sky130_fd_sc_hd__nor2_2
Xinput208 W1END[2] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_4
Xinput219 W2MID[1] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1087_ Inst_RegFile_32x4/_0452_ Inst_RegFile_32x4/_0453_ Inst_RegFile_32x4/_0454_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0513_ sky130_fd_sc_hd__or3b_4
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2 net226
+ AD0 AD1 AD2 ConfigBits\[362\] ConfigBits\[363\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame10_bit27 net68 net82 VGND VGND VPWR VPWR ConfigBits\[89\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit16 net56 net82 VGND VGND VPWR VPWR ConfigBits\[78\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame6_bit30 net72 net97 VGND VGND VPWR VPWR ConfigBits\[220\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_31__0_ FrameData_O_i\[31\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__1010_ Inst_RegFile_32x4/_0451_ Inst_RegFile_32x4__1340_/Q Inst_RegFile_32x4/_0459_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0725_ Inst_RegFile_32x4/_0151_ Inst_RegFile_32x4/_0164_ Inst_RegFile_32x4/_0181_
+ Inst_RegFile_32x4/_0190_ A_ADR3 A_ADR4 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0191_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1 net11
+ net155 net163 net206 ConfigBits\[274\] ConfigBits\[275\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xdata_outbuf_22__0_ FrameData_O_i\[22\] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1208_ Inst_RegFile_32x4/_0458_ Inst_RegFile_32x4/_0571_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0586_ sky130_fd_sc_hd__nand2_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG1 net129 net197 net212 JE2BEG\[4\]
+ ConfigBits\[408\] ConfigBits\[409\] VGND VGND VPWR VPWR J_l_GH_BEG\[1\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1139_ Inst_RegFile_32x4/_0451_ Inst_RegFile_32x4__1392_/Q Inst_RegFile_32x4/_0544_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_outbuf_13__0_ FrameData_O_i\[13\] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame9_bit23 net64 net100 VGND VGND VPWR VPWR ConfigBits\[117\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit12 net52 net100 VGND VGND VPWR VPWR ConfigBits\[106\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame5_bit9 net80 net96 VGND VGND VPWR VPWR ConfigBits\[231\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XS4BEG_outbuf_2__0_ S4BEG_i\[2\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix__60_ net222 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst1 BD1 J2MID_ABb_BEG\[1\]
+ J2MID_CDb_BEG\[1\] J2END_GH_BEG\[3\] ConfigBits\[74\] ConfigBits\[75\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0 net101
+ net105 net1 net5 ConfigBits\[314\] ConfigBits\[315\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2 net229
+ AD0 AD1 AD3 ConfigBits\[326\] ConfigBits\[327\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0708_ Inst_RegFile_32x4/_0130_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0174_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2 BD0 BD1
+ BD2 BD3 ConfigBits\[106\] ConfigBits\[107\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XS4END_inbuf_0__0_ net183 VGND VGND VPWR VPWR S4BEG_i\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_54_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput309 net309 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0990_ Inst_RegFile_32x4__1427_/Q Inst_RegFile_32x4__1423_/Q Inst_RegFile_32x4/_0326_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1473_ net205 Inst_RegFile_32x4/_0125_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1473_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XNN4END_inbuf_8__0_ net140 VGND VGND VPWR VPWR NN4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_2
XEE4BEG_outbuf_1__0_ EE4BEG_i\[1\] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_1
XW6END_inbuf_4__0_ net234 VGND VGND VPWR VPWR W6BEG_i\[4\] sky130_fd_sc_hd__clkbuf_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__43_ net168 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame12_bit19 net59 net84 VGND VGND VPWR VPWR ConfigBits\[17\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit11 net51 net99 VGND VGND VPWR VPWR ConfigBits\[137\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit22 net63 net99 VGND VGND VPWR VPWR ConfigBits\[148\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG0 net119 net19 net224
+ JN2BEG\[5\] ConfigBits\[174\] ConfigBits\[175\] VGND VGND VPWR VPWR J2MID_EFa_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[290\] ConfigBits\[291\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame12_bit8 net79 net84 VGND VGND VPWR VPWR ConfigBits\[6\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0973_ Inst_RegFile_32x4/_0306_ Inst_RegFile_32x4/_0424_ Inst_RegFile_32x4/_0340_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1456_ net205 Inst_RegFile_32x4/_0108_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1456_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__1_/A1 ConfigBits\[76\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix__26_ net115 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1387_ net205 Inst_RegFile_32x4__1387_/D VGND VGND VPWR VPWR Inst_RegFile_32x4__1387_/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 E2MID[6] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame1_bit1 net60 net92 VGND VGND VPWR VPWR ConfigBits\[351\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG1 net116 net16 net168
+ net221 ConfigBits\[216\] ConfigBits\[217\] VGND VGND VPWR VPWR J2MID_GHb_BEG\[1\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame11_bit18 net58 net83 VGND VGND VPWR VPWR ConfigBits\[48\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1310_ Inst_RegFile_32x4/_0645_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0114_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame11_bit29 net70 net83 VGND VGND VPWR VPWR ConfigBits\[59\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1241_ Inst_RegFile_32x4/_0577_ Inst_RegFile_32x4__1432_/Q Inst_RegFile_32x4/_0606_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0607_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1172_ Inst_RegFile_32x4/_0563_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0058_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame7_bit10 net50 net98 VGND VGND VPWR VPWR ConfigBits\[168\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame7_bit21 net62 net98 VGND VGND VPWR VPWR ConfigBits\[179\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0956_ Inst_RegFile_32x4__1426_/Q Inst_RegFile_32x4__1422_/Q Inst_RegFile_32x4/_0326_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0410_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0887_ Inst_RegFile_32x4/_0343_ Inst_RegFile_32x4/_0344_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0345_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG3 net105 net40 net157 net210
+ ConfigBits\[236\] ConfigBits\[237\] VGND VGND VPWR VPWR J2END_CD_BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1439_ net205 Inst_RegFile_32x4/_0091_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1439_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput470 net470 VGND VGND VPWR VPWR W2BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix__09_ net14 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__buf_1
Xoutput481 net481 VGND VGND VPWR VPWR W6BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput492 net492 VGND VGND VPWR VPWR WW4BEG[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XEE4BEG_outbuf_11__0_ EE4BEG_i\[11\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_cus_mux41_buf_inst0 net108 net160
+ J2MID_CDa_BEG\[1\] J2MID_CDb_BEG\[2\] ConfigBits\[155\] ConfigBits\[156\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame8_bit7 net78 net99 VGND VGND VPWR VPWR ConfigBits\[133\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0810_ Inst_RegFile_32x4__1443_/Q Inst_RegFile_32x4__1439_/Q Inst_RegFile_32x4/_0174_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0672_ Inst_RegFile_32x4__1404_/Q Inst_RegFile_32x4__1380_/Q Inst_RegFile_32x4/_0137_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0741_ Inst_RegFile_32x4/_0202_ Inst_RegFile_32x4/_0204_ Inst_RegFile_32x4/_0205_
+ Inst_RegFile_32x4/_0149_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0206_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__1224_ D2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0596_ sky130_fd_sc_hd__clkbuf_2
Xinput209 W1END[3] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_4
XInst_RegFile_32x4__1086_ Inst_RegFile_32x4/_0512_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0023_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1155_ Inst_RegFile_32x4/_0553_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0051_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0939_ Inst_RegFile_32x4/_0306_ Inst_RegFile_32x4/_0392_ Inst_RegFile_32x4/_0340_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0393_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[362\] ConfigBits\[363\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_outbuf_0__0_ FrameData_O_i\[0\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame10_bit28 net69 net82 VGND VGND VPWR VPWR ConfigBits\[90\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit17 net57 net82 VGND VGND VPWR VPWR ConfigBits\[79\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame6_bit20 net61 net97 VGND VGND VPWR VPWR ConfigBits\[210\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit31 net73 net97 VGND VGND VPWR VPWR ConfigBits\[221\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_inbuf_24__0_ net65 VGND VGND VPWR VPWR FrameData_O_i\[24\] sky130_fd_sc_hd__buf_1
XFILLER_0_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0724_ Inst_RegFile_32x4/_0184_ Inst_RegFile_32x4/_0187_ Inst_RegFile_32x4/_0189_
+ Inst_RegFile_32x4/_0163_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0190_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2 net208
+ AD0 AD1 AD2 ConfigBits\[274\] ConfigBits\[275\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1207_ Inst_RegFile_32x4/_0585_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0071_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_3__0_ net94 VGND VGND VPWR VPWR FrameStrobe_O_i\[3\] sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_15__0_ net55 VGND VGND VPWR VPWR FrameData_O_i\[15\] sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__1069_ Inst_RegFile_32x4/_0473_ Inst_RegFile_32x4/_0502_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0503_ sky130_fd_sc_hd__nor2_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG2 net24 net180 net247 JS2BEG\[4\]
+ ConfigBits\[410\] ConfigBits\[411\] VGND VGND VPWR VPWR J_l_GH_BEG\[2\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1138_ Inst_RegFile_32x4/_0458_ Inst_RegFile_32x4/_0471_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0544_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame9_bit13 net53 net100 VGND VGND VPWR VPWR ConfigBits\[107\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit24 net65 net100 VGND VGND VPWR VPWR ConfigBits\[118\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1 net33
+ net153 net155 net157 ConfigBits\[314\] ConfigBits\[315\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[326\] ConfigBits\[327\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0707_ Inst_RegFile_32x4/_0128_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0173_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3 J2MID_ABb_BEG\[1\]
+ J2MID_CDb_BEG\[1\] J2MID_EFb_BEG\[1\] J2MID_GHb_BEG\[1\] ConfigBits\[106\] ConfigBits\[107\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame5_bit30 net72 net96 VGND VGND VPWR VPWR ConfigBits\[252\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_outbuf_18__0_ FrameStrobe_O_i\[18\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1472_ net205 Inst_RegFile_32x4/_0124_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1472_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__42_ net167 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkbuf_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG0 net146 net182 net238 JN2BEG\[1\]
+ ConfigBits\[382\] ConfigBits\[383\] VGND VGND VPWR VPWR J_l_AB_BEG\[0\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame8_bit12 net52 net99 VGND VGND VPWR VPWR ConfigBits\[138\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit23 net64 net99 VGND VGND VPWR VPWR ConfigBits\[149\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XWW4END_inbuf_9__0_ net242 VGND VGND VPWR VPWR WW4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG1 net115 net15 net167
+ JE2BEG\[5\] ConfigBits\[176\] ConfigBits\[177\] VGND VGND VPWR VPWR J2MID_EFa_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3/X ConfigBits\[292\]
+ ConfigBits\[293\] VGND VGND VPWR VPWR JE2BEG\[1\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame12_bit9 net80 net84 VGND VGND VPWR VPWR ConfigBits\[7\]
+ Inst_RegFile_ConfigMem_Inst_frame12_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0972_ Inst_RegFile_32x4__1371_/Q Inst_RegFile_32x4__1367_/Q Inst_RegFile_32x4/_0338_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1455_ net205 Inst_RegFile_32x4/_0107_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1455_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1386_ net205 Inst_RegFile_32x4__1386_/D VGND VGND VPWR VPWR Inst_RegFile_32x4__1386_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__25_ net114 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame1_bit2 net71 net92 VGND VGND VPWR VPWR ConfigBits\[352\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG2 net118 net18 net170
+ net223 ConfigBits\[218\] ConfigBits\[219\] VGND VGND VPWR VPWR J2MID_GHb_BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
Xstrobe_outbuf_0__0_ FrameStrobe_O_i\[0\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1240_ Inst_RegFile_32x4/_0554_ Inst_RegFile_32x4/_0600_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0606_ sky130_fd_sc_hd__nand2_2
XInst_RegFile_ConfigMem_Inst_frame11_bit19 net59 net83 VGND VGND VPWR VPWR ConfigBits\[49\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1171_ Inst_RegFile_32x4__1406_/Q Inst_RegFile_32x4/_0530_ Inst_RegFile_32x4/_0560_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0563_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame7_bit11 net51 net98 VGND VGND VPWR VPWR ConfigBits\[169\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame7_bit22 net63 net98 VGND VGND VPWR VPWR ConfigBits\[180\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0955_ Inst_RegFile_32x4/_0402_ Inst_RegFile_32x4/_0404_ Inst_RegFile_32x4/_0406_
+ Inst_RegFile_32x4/_0408_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0409_ sky130_fd_sc_hd__o22a_2
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0886_ Inst_RegFile_32x4__1424_/Q Inst_RegFile_32x4__1420_/Q Inst_RegFile_32x4/_0292_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0344_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1438_ net205 Inst_RegFile_32x4/_0090_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1438_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1369_ net205 Inst_RegFile_32x4/_0029_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1369_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput482 net482 VGND VGND VPWR VPWR W6BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput493 net493 VGND VGND VPWR VPWR WW4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput460 net460 VGND VGND VPWR VPWR W1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput471 net471 VGND VGND VPWR VPWR W2BEGb[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix__08_ net13 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__buf_1
XFILLER_0_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_15__0_ net87 VGND VGND VPWR VPWR FrameStrobe_O_i\[15\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_cus_mux41_buf_inst1 J2END_GH_BEG\[3\]
+ JN2BEG\[0\] JS2BEG\[0\] JW2BEG\[0\] ConfigBits\[155\] ConfigBits\[156\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_en_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XE6END_inbuf_9__0_ net23 VGND VGND VPWR VPWR E6BEG_i\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame8_bit8 net79 net99 VGND VGND VPWR VPWR ConfigBits\[134\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0671_ Inst_RegFile_32x4/_0136_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0137_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0740_ Inst_RegFile_32x4__1345_/Q Inst_RegFile_32x4__1393_/Q Inst_RegFile_32x4__1465_/Q
+ Inst_RegFile_32x4__1461_/Q Inst_RegFile_32x4/_0146_ Inst_RegFile_32x4/_0161_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0205_ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1223_ Inst_RegFile_32x4/_0595_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0077_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1085_ Inst_RegFile_32x4__1363_/Q Inst_RegFile_32x4/_0500_ Inst_RegFile_32x4/_0508_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0512_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1154_ Inst_RegFile_32x4__1399_/Q Inst_RegFile_32x4/_0532_ Inst_RegFile_32x4/_0549_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0553_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0938_ Inst_RegFile_32x4__1370_/Q Inst_RegFile_32x4__1366_/Q Inst_RegFile_32x4/_0338_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0392_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0869_ Inst_RegFile_32x4__1456_/Q Inst_RegFile_32x4__1452_/Q Inst_RegFile_32x4/_0326_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3/X ConfigBits\[364\]
+ ConfigBits\[365\] VGND VGND VPWR VPWR JW2BEG\[3\] sky130_fd_sc_hd__mux4_2
Xoutput290 net290 VGND VGND VPWR VPWR EE4BEG[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XE6BEG_outbuf_1__0_ E6BEG_i\[1\] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame10_bit18 net58 net82 VGND VGND VPWR VPWR ConfigBits\[80\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame10_bit29 net70 net82 VGND VGND VPWR VPWR ConfigBits\[91\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame6_bit21 net62 net97 VGND VGND VPWR VPWR ConfigBits\[211\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit10 net50 net97 VGND VGND VPWR VPWR ConfigBits\[200\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XN4END_inbuf_0__0_ net131 VGND VGND VPWR VPWR N4BEG_i\[0\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0723_ Inst_RegFile_32x4__1408_/Q Inst_RegFile_32x4__1340_/Q Inst_RegFile_32x4__1400_/Q
+ Inst_RegFile_32x4__1468_/Q Inst_RegFile_32x4/_0160_ Inst_RegFile_32x4/_0188_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0189_ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3 AD3 BD0
+ BD2 BD3 ConfigBits\[274\] ConfigBits\[275\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1206_ Inst_RegFile_32x4/_0584_ Inst_RegFile_32x4__1419_/Q Inst_RegFile_32x4/_0578_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0585_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1137_ Inst_RegFile_32x4/_0543_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0043_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1068_ Inst_RegFile_32x4/_0452_ Inst_RegFile_32x4/_0453_ Inst_RegFile_32x4/_0454_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0502_ sky130_fd_sc_hd__or3_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG3 net137 net21 net210 JW2BEG\[4\]
+ ConfigBits\[412\] ConfigBits\[413\] VGND VGND VPWR VPWR J_l_GH_BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_66_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame9_bit14 net54 net100 VGND VGND VPWR VPWR ConfigBits\[108\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit25 net66 net100 VGND VGND VPWR VPWR ConfigBits\[119\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_7__0_ net78 VGND VGND VPWR VPWR FrameData_O_i\[7\] sky130_fd_sc_hd__buf_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__0706_ Inst_RegFile_32x4/_0168_ Inst_RegFile_32x4/_0170_ Inst_RegFile_32x4/_0171_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0172_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2 net206
+ AD0 AD1 AD2 ConfigBits\[314\] ConfigBits\[315\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3/X ConfigBits\[328\]
+ ConfigBits\[329\] VGND VGND VPWR VPWR JS2BEG\[2\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3/X ConfigBits\[108\]
+ ConfigBits\[109\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame5_bit20 net61 net96 VGND VGND VPWR VPWR ConfigBits\[242\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame5_bit31 net73 net96 VGND VGND VPWR VPWR ConfigBits\[253\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame4_bit0 net49 net95 VGND VGND VPWR VPWR ConfigBits\[254\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1471_ net205 Inst_RegFile_32x4/_0123_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1471_/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__41_ net166 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkbuf_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG1 net41 net181 net217 JE2BEG\[1\]
+ ConfigBits\[384\] ConfigBits\[385\] VGND VGND VPWR VPWR J_l_AB_BEG\[1\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame8_bit13 net53 net99 VGND VGND VPWR VPWR ConfigBits\[139\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame8_bit24 net65 net99 VGND VGND VPWR VPWR ConfigBits\[150\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG2 net117 net169 net222
+ JS2BEG\[5\] ConfigBits\[178\] ConfigBits\[179\] VGND VGND VPWR VPWR J2MID_EFa_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput190 SS4END[10] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
XNN4BEG_outbuf_1__0_ NN4BEG_i\[1\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0971_ Inst_RegFile_32x4/_0334_ Inst_RegFile_32x4/_0422_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0423_ sky130_fd_sc_hd__and2b_1
XN4BEG_outbuf_5__0_ N4BEG_i\[5\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame4_bit30 net72 net95 VGND VGND VPWR VPWR ConfigBits\[284\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1454_ net205 Inst_RegFile_32x4/_0106_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1454_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1385_ net205 Inst_RegFile_32x4__1385_/D VGND VGND VPWR VPWR Inst_RegFile_32x4__1385_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__24_ net113 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSS4BEG_outbuf_4__0_ SS4BEG_i\[4\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame1_bit3 net74 net92 VGND VGND VPWR VPWR ConfigBits\[353\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG3 net114 net14 net166
+ net219 ConfigBits\[220\] ConfigBits\[221\] VGND VGND VPWR VPWR J2MID_GHb_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1170_ Inst_RegFile_32x4/_0562_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0057_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XW6BEG_outbuf_5__0_ W6BEG_i\[5\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame7_bit23 net64 net98 VGND VGND VPWR VPWR ConfigBits\[181\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame7_bit12 net52 net98 VGND VGND VPWR VPWR ConfigBits\[170\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0954_ Inst_RegFile_32x4/_0296_ Inst_RegFile_32x4/_0407_ Inst_RegFile_32x4/_0340_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0408_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0885_ Inst_RegFile_32x4/_0289_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0343_
+ sky130_fd_sc_hd__buf_1
XFILLER_0_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1299_ Inst_RegFile_32x4/_0639_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0109_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1437_ net205 Inst_RegFile_32x4/_0089_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1437_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1368_ net205 Inst_RegFile_32x4/_0028_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1368_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput494 net494 VGND VGND VPWR VPWR WW4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput483 net483 VGND VGND VPWR VPWR W6BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput450 net450 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput461 net461 VGND VGND VPWR VPWR W1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput472 net472 VGND VGND VPWR VPWR W2BEGb[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix__07_ JE2BEG\[7\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0 net106
+ net128 net4 net6 ConfigBits\[254\] ConfigBits\[255\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame8_bit9 net80 net99 VGND VGND VPWR VPWR ConfigBits\[135\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_D0 J2MID_ABa_BEG\[0\] J2MID_ABb_BEG\[0\]
+ J2END_AB_BEG\[0\] J_l_AB_BEG\[0\] ConfigBits\[136\] ConfigBits\[137\] VGND VGND
+ VPWR VPWR D0 sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__0670_ A_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0136_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1222_ Inst_RegFile_32x4__1425_/Q Inst_RegFile_32x4/_0594_ Inst_RegFile_32x4/_0592_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0595_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1153_ Inst_RegFile_32x4/_0552_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0050_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1084_ Inst_RegFile_32x4/_0511_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0022_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0868_ B_ADR0 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0326_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0937_ Inst_RegFile_32x4/_0334_ Inst_RegFile_32x4/_0390_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0391_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_outbuf_25__0_ FrameData_O_i\[25\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0799_ Inst_RegFile_32x4/_0255_ Inst_RegFile_32x4/_0257_ Inst_RegFile_32x4/_0259_
+ Inst_RegFile_32x4/_0261_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0262_ sky130_fd_sc_hd__o22a_1
Xoutput280 net280 VGND VGND VPWR VPWR E6BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput291 net291 VGND VGND VPWR VPWR EE4BEG[14] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_ConfigMem_Inst_frame10_bit19 net59 net82 VGND VGND VPWR VPWR ConfigBits\[81\]
+ Inst_RegFile_ConfigMem_Inst_frame10_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit11 net51 net97 VGND VGND VPWR VPWR ConfigBits\[201\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit22 net63 net97 VGND VGND VPWR VPWR ConfigBits\[212\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_16__0_ FrameData_O_i\[16\] VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XS4BEG_outbuf_5__0_ S4BEG_i\[5\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0722_ A_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0188_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3/X ConfigBits\[276\]
+ ConfigBits\[277\] VGND VGND VPWR VPWR JN2BEG\[5\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__1205_ Inst_RegFile_32x4/_0467_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0584_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_32x4__1136_ Inst_RegFile_32x4__1383_/Q Inst_RegFile_32x4/_0532_ Inst_RegFile_32x4/_0539_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0543_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1067_ Inst_RegFile_32x4/_0501_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0015_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame9_bit15 net55 net100 VGND VGND VPWR VPWR ConfigBits\[109\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit26 net67 net100 VGND VGND VPWR VPWR ConfigBits\[120\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XS4END_inbuf_3__0_ net186 VGND VGND VPWR VPWR S4BEG_i\[3\] sky130_fd_sc_hd__buf_2
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0705_ A_ADR2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0171_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3 AD3 BD0
+ BD1 BD2 ConfigBits\[314\] ConfigBits\[315\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XEE4BEG_outbuf_4__0_ EE4BEG_i\[4\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XW6END_inbuf_7__0_ net237 VGND VGND VPWR VPWR W6BEG_i\[7\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame5_bit21 net62 net96 VGND VGND VPWR VPWR ConfigBits\[243\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1119_ Inst_RegFile_32x4/_0533_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0035_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame5_bit10 net50 net96 VGND VGND VPWR VPWR ConfigBits\[232\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame4_bit1 net60 net95 VGND VGND VPWR VPWR ConfigBits\[255\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1470_ net205 Inst_RegFile_32x4/_0122_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1470_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix__40_ net165 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit14 net54 net99 VGND VGND VPWR VPWR ConfigBits\[140\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG2 net128 net24 net229 JS2BEG\[1\]
+ ConfigBits\[386\] ConfigBits\[387\] VGND VGND VPWR VPWR J_l_AB_BEG\[2\] sky130_fd_sc_hd__mux4_1
XFILLER_0_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame8_bit25 net66 net99 VGND VGND VPWR VPWR ConfigBits\[151\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG3 net13 net165 net218
+ JW2BEG\[5\] ConfigBits\[180\] ConfigBits\[181\] VGND VGND VPWR VPWR J2MID_EFa_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput180 S4END[1] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_4
Xinput191 SS4END[11] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0970_ Inst_RegFile_32x4__1379_/Q Inst_RegFile_32x4__1375_/Q Inst_RegFile_32x4/_0335_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0422_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame4_bit20 net61 net95 VGND VGND VPWR VPWR ConfigBits\[274\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1453_ net205 Inst_RegFile_32x4/_0105_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1453_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_ConfigMem_Inst_frame4_bit31 net73 net95 VGND VGND VPWR VPWR ConfigBits\[285\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix__23_ JN2BEG\[7\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1384_ net205 Inst_RegFile_32x4__1384_/D VGND VGND VPWR VPWR Inst_RegFile_32x4__1384_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_S1BEG0 BD0 J2MID_CDb_BEG\[3\] JE2BEG\[3\]
+ J_l_CD_BEG\[1\] ConfigBits\[58\] ConfigBits\[59\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__mux4_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame1_bit4 net75 net92 VGND VGND VPWR VPWR ConfigBits\[354\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame11_bit0 net49 net83 VGND VGND VPWR VPWR ConfigBits\[30\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame7_bit24 net65 net98 VGND VGND VPWR VPWR ConfigBits\[182\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame7_bit13 net53 net98 VGND VGND VPWR VPWR ConfigBits\[171\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0953_ Inst_RegFile_32x4__1434_/Q Inst_RegFile_32x4__1430_/Q Inst_RegFile_32x4/_0338_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0407_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0884_ Inst_RegFile_32x4/_0328_ Inst_RegFile_32x4/_0333_ Inst_RegFile_32x4/_0337_
+ Inst_RegFile_32x4/_0341_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0342_ sky130_fd_sc_hd__o22a_1
XN4END_inbuf_11__0_ net127 VGND VGND VPWR VPWR N4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1436_ net205 Inst_RegFile_32x4/_0088_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1436_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4END_inbuf_10__0_ net194 VGND VGND VPWR VPWR SS4BEG_i\[10\] sky130_fd_sc_hd__buf_2
XInst_RegFile_32x4__1298_ Inst_RegFile_32x4__1457_/Q Inst_RegFile_32x4/_0461_ Inst_RegFile_32x4/_0637_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0639_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1367_ net205 Inst_RegFile_32x4/_0027_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1367_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_switch_matrix__06_ JE2BEG\[6\] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_1
Xoutput484 net484 VGND VGND VPWR VPWR W6BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput495 net495 VGND VGND VPWR VPWR WW4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput451 net451 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput440 net440 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput462 net462 VGND VGND VPWR VPWR W1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput473 net473 VGND VGND VPWR VPWR W2BEGb[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_3__0_ FrameData_O_i\[3\] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1 net33
+ net24 net158 net211 ConfigBits\[254\] ConfigBits\[255\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame3_bit30 net72 net94 VGND VGND VPWR VPWR ConfigBits\[316\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_D1 J2MID_ABa_BEG\[1\] J2MID_ABb_BEG\[1\]
+ J2END_AB_BEG\[1\] J_l_AB_BEG\[1\] ConfigBits\[138\] ConfigBits\[139\] VGND VGND
+ VPWR VPWR D1 sky130_fd_sc_hd__mux4_2
XFILLER_0_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1221_ D1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0594_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1152_ Inst_RegFile_32x4__1398_/Q Inst_RegFile_32x4/_0530_ Inst_RegFile_32x4/_0549_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1083_ Inst_RegFile_32x4__1362_/Q Inst_RegFile_32x4/_0498_ Inst_RegFile_32x4/_0508_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_27__0_ net68 VGND VGND VPWR VPWR FrameData_O_i\[27\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0798_ Inst_RegFile_32x4/_0145_ Inst_RegFile_32x4/_0260_ Inst_RegFile_32x4/_0179_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0261_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0936_ Inst_RegFile_32x4__1378_/Q Inst_RegFile_32x4__1374_/Q Inst_RegFile_32x4/_0303_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0867_ Inst_RegFile_32x4/_0316_ Inst_RegFile_32x4/_0320_ Inst_RegFile_32x4/_0323_
+ Inst_RegFile_32x4/_0324_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0325_ sky130_fd_sc_hd__o22a_1
XInst_RegFile_32x4__1419_ net205 Inst_RegFile_32x4/_0071_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1419_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput270 net270 VGND VGND VPWR VPWR E2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xstrobe_inbuf_6__0_ net97 VGND VGND VPWR VPWR FrameStrobe_O_i\[6\] sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_18__0_ net58 VGND VGND VPWR VPWR FrameData_O_i\[18\] sky130_fd_sc_hd__clkbuf_1
Xoutput281 net281 VGND VGND VPWR VPWR E6BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput292 net292 VGND VGND VPWR VPWR EE4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0 net102
+ net108 net130 net8 ConfigBits\[294\] ConfigBits\[295\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame6_bit12 net52 net97 VGND VGND VPWR VPWR ConfigBits\[202\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame6_bit23 net64 net97 VGND VGND VPWR VPWR ConfigBits\[213\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0721_ Inst_RegFile_32x4/_0185_ Inst_RegFile_32x4/_0186_ Inst_RegFile_32x4/_0139_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0187_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1204_ Inst_RegFile_32x4/_0583_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0070_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1135_ Inst_RegFile_32x4/_0542_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0042_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1066_ Inst_RegFile_32x4__1355_/Q Inst_RegFile_32x4/_0500_ Inst_RegFile_32x4/_0494_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0919_ Inst_RegFile_32x4__1433_/Q Inst_RegFile_32x4__1429_/Q Inst_RegFile_32x4/_0338_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0375_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame9_bit16 net56 net100 VGND VGND VPWR VPWR ConfigBits\[110\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame9_bit27 net68 net100 VGND VGND VPWR VPWR ConfigBits\[121\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XS4END_inbuf_11__0_ net179 VGND VGND VPWR VPWR S4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3/X ConfigBits\[316\]
+ ConfigBits\[317\] VGND VGND VPWR VPWR JE2BEG\[7\] sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__0704_ Inst_RegFile_32x4__1448_/Q Inst_RegFile_32x4__1472_/Q Inst_RegFile_32x4/_0169_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst0 net104
+ net4 net209 AD2 ConfigBits\[21\] ConfigBits\[22\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1118_ Inst_RegFile_32x4__1375_/Q Inst_RegFile_32x4/_0532_ Inst_RegFile_32x4/_0526_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0533_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame5_bit11 net51 net96 VGND VGND VPWR VPWR ConfigBits\[233\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame5_bit22 net63 net96 VGND VGND VPWR VPWR ConfigBits\[244\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1049_ Inst_RegFile_32x4__1350_/Q Inst_RegFile_32x4/_0479_ Inst_RegFile_32x4/_0486_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame4_bit2 net71 net95 VGND VGND VPWR VPWR ConfigBits\[256\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0 net102
+ net110 net2 net10 ConfigBits\[366\] ConfigBits\[367\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame8_bit26 net67 net99 VGND VGND VPWR VPWR ConfigBits\[152\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit15 net55 net99 VGND VGND VPWR VPWR ConfigBits\[141\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSS4END_inbuf_1__0_ net200 VGND VGND VPWR VPWR SS4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_2
XEE4END_inbuf_10__0_ net38 VGND VGND VPWR VPWR EE4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG3 net121 net21 net173 JW2BEG\[1\]
+ ConfigBits\[388\] ConfigBits\[389\] VGND VGND VPWR VPWR J_l_AB_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_35_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput192 SS4END[12] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
Xinput181 S4END[2] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xinput170 S2MID[5] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_2
XFILLER_0_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xstrobe_outbuf_3__0_ FrameStrobe_O_i\[3\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame4_bit21 net62 net95 VGND VGND VPWR VPWR ConfigBits\[275\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1452_ net205 Inst_RegFile_32x4/_0104_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1452_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_ConfigMem_Inst_frame4_bit10 net50 net95 VGND VGND VPWR VPWR ConfigBits\[264\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix__22_ JN2BEG\[6\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1383_ net205 Inst_RegFile_32x4/_0043_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1383_/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_S1BEG1 BD1 J2MID_EFb_BEG\[0\] JE2BEG\[0\]
+ J_l_EF_BEG\[2\] ConfigBits\[60\] ConfigBits\[61\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__mux4_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame1_bit5 net76 net92 VGND VGND VPWR VPWR ConfigBits\[355\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XEE4END_inbuf_0__0_ net43 VGND VGND VPWR VPWR EE4BEG_i\[0\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame11_bit1 net60 net83 VGND VGND VPWR VPWR ConfigBits\[31\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XWW4BEG_outbuf_1__0_ WW4BEG_i\[1\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_18__0_ net90 VGND VGND VPWR VPWR FrameStrobe_O_i\[18\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame7_bit25 net66 net98 VGND VGND VPWR VPWR ConfigBits\[183\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_B_ADR0 J2MID_GHa_BEG\[0\] J2MID_GHb_BEG\[0\]
+ J2END_GH_BEG\[0\] J_l_GH_BEG\[0\] ConfigBits\[125\] ConfigBits\[126\] VGND VGND
+ VPWR VPWR B_ADR0 sky130_fd_sc_hd__mux4_2
XFILLER_0_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame7_bit14 net54 net98 VGND VGND VPWR VPWR ConfigBits\[172\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0952_ Inst_RegFile_32x4/_0290_ Inst_RegFile_32x4/_0405_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0406_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_cus_mux41_buf_inst0 net106 net158
+ J2MID_GHa_BEG\[1\] J2MID_GHb_BEG\[2\] ConfigBits\[122\] ConfigBits\[123\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0 net145
+ net3 net197 net208 ConfigBits\[110\] ConfigBits\[111\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0 net109
+ net3 net9 net42 ConfigBits\[330\] ConfigBits\[331\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0883_ Inst_RegFile_32x4/_0306_ Inst_RegFile_32x4/_0339_ Inst_RegFile_32x4/_0340_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0341_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1435_ net205 Inst_RegFile_32x4/_0087_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1435_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1366_ net205 Inst_RegFile_32x4/_0026_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1366_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput452 net452 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput430 net430 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput441 net441 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1297_ Inst_RegFile_32x4/_0638_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0108_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix__05_ JE2BEG\[5\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_1
Xoutput485 net485 VGND VGND VPWR VPWR W6BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput496 net496 VGND VGND VPWR VPWR WW4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput463 net463 VGND VGND VPWR VPWR W2BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput474 net474 VGND VGND VPWR VPWR W2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XE6BEG_outbuf_4__0_ E6BEG_i\[4\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG0 net120 net20 net172
+ net225 ConfigBits\[190\] ConfigBits\[191\] VGND VGND VPWR VPWR J2MID_ABb_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2 net229
+ AD1 AD2 AD3 ConfigBits\[254\] ConfigBits\[255\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame3_bit20 net61 net94 VGND VGND VPWR VPWR ConfigBits\[306\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit31 net73 net94 VGND VGND VPWR VPWR ConfigBits\[317\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_D2 J2MID_ABa_BEG\[2\] J2MID_ABb_BEG\[2\]
+ J2END_AB_BEG\[2\] J_l_AB_BEG\[2\] ConfigBits\[140\] ConfigBits\[141\] VGND VGND
+ VPWR VPWR D2 sky130_fd_sc_hd__mux4_2
XInst_RegFile_32x4__1220_ Inst_RegFile_32x4/_0593_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0076_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__1151_ Inst_RegFile_32x4/_0551_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0049_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1082_ Inst_RegFile_32x4/_0510_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0021_
+ sky130_fd_sc_hd__clkbuf_1
XN4END_inbuf_3__0_ net134 VGND VGND VPWR VPWR N4BEG_i\[3\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__0935_ Inst_RegFile_32x4/_0346_ Inst_RegFile_32x4/_0388_ Inst_RegFile_32x4/_0300_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0797_ Inst_RegFile_32x4__1371_/Q Inst_RegFile_32x4__1367_/Q Inst_RegFile_32x4/_0177_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0866_ Inst_RegFile_32x4/_0309_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0324_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1418_ net205 Inst_RegFile_32x4/_0070_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1418_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput282 net282 VGND VGND VPWR VPWR E6BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput293 net293 VGND VGND VPWR VPWR EE4BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput271 net271 VGND VGND VPWR VPWR E2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput260 net260 VGND VGND VPWR VPWR E2BEG[2] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1349_ net205 Inst_RegFile_32x4/_0009_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1349_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_ConfigMem_Inst_frame7_bit0 net49 net98 VGND VGND VPWR VPWR ConfigBits\[158\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1 net24
+ net160 net197 net213 ConfigBits\[294\] ConfigBits\[295\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame6_bit13 net53 net97 VGND VGND VPWR VPWR ConfigBits\[203\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit24 net65 net97 VGND VGND VPWR VPWR ConfigBits\[214\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__0720_ Inst_RegFile_32x4__1416_/Q Inst_RegFile_32x4__1412_/Q Inst_RegFile_32x4/_0169_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0186_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1203_ Inst_RegFile_32x4/_0582_ Inst_RegFile_32x4__1418_/Q Inst_RegFile_32x4/_0578_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0583_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1065_ Inst_RegFile_32x4/_0467_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0500_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1134_ Inst_RegFile_32x4__1382_/Q Inst_RegFile_32x4/_0530_ Inst_RegFile_32x4/_0539_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0542_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0918_ Inst_RegFile_32x4/_0334_ Inst_RegFile_32x4/_0373_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0374_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_ConfigMem_Inst_frame2_bit30 net72 net93 VGND VGND VPWR VPWR ConfigBits\[348\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0849_ Inst_RegFile_32x4/_0297_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0307_
+ sky130_fd_sc_hd__buf_2
XInst_RegFile_ConfigMem_Inst_frame9_bit28 net69 net100 VGND VGND VPWR VPWR ConfigBits\[122\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit17 net57 net100 VGND VGND VPWR VPWR ConfigBits\[111\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0703_ Inst_RegFile_32x4/_0130_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0169_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst1 BD2 J2MID_ABa_BEG\[2\]
+ J2MID_CDa_BEG\[2\] J2END_EF_BEG\[1\] ConfigBits\[21\] ConfigBits\[22\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1117_ D3 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0532_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame5_bit12 net52 net96 VGND VGND VPWR VPWR ConfigBits\[234\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1048_ Inst_RegFile_32x4/_0488_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0009_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame5_bit23 net64 net96 VGND VGND VPWR VPWR ConfigBits\[245\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst0 net102
+ net154 net207 AD0 ConfigBits\[103\] ConfigBits\[104\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame4_bit3 net74 net95 VGND VGND VPWR VPWR ConfigBits\[257\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 J2MID_EFb_BEG\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1 net154
+ net156 net162 net207 ConfigBits\[366\] ConfigBits\[367\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XN4BEG_outbuf_8__0_ N4BEG_i\[8\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_1
XNN4BEG_outbuf_4__0_ NN4BEG_i\[4\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkbuf_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit27 net68 net99 VGND VGND VPWR VPWR ConfigBits\[153\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame8_bit16 net56 net99 VGND VGND VPWR VPWR ConfigBits\[142\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSS4BEG_outbuf_7__0_ SS4BEG_i\[7\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4BEG_outbuf_11__0_ S4BEG_i\[11\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput193 SS4END[13] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
Xinput182 S4END[3] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_2
Xinput171 S2MID[6] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
Xinput160 S2END[3] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0 net104
+ net112 net144 net4 ConfigBits\[278\] ConfigBits\[279\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame4_bit22 net63 net95 VGND VGND VPWR VPWR ConfigBits\[276\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1451_ net205 Inst_RegFile_32x4/_0103_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1451_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_ConfigMem_Inst_frame4_bit11 net51 net95 VGND VGND VPWR VPWR ConfigBits\[265\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1382_ net205 Inst_RegFile_32x4/_0042_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1382_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix__21_ JN2BEG\[5\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
XW6BEG_outbuf_8__0_ W6BEG_i\[8\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__clkbuf_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_S1BEG2 BD2 J2MID_GHb_BEG\[1\] JE2BEG\[1\]
+ J_l_GH_BEG\[3\] ConfigBits\[62\] ConfigBits\[63\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__mux4_1
XFILLER_0_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame1_bit6 net77 net92 VGND VGND VPWR VPWR ConfigBits\[356\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame11_bit2 net71 net83 VGND VGND VPWR VPWR ConfigBits\[32\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__1_/A1 ConfigBits\[49\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst0 net104
+ net4 net209 AD2 ConfigBits\[77\] ConfigBits\[78\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__1_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_B_ADR1 J2MID_GHa_BEG\[1\] J2MID_GHb_BEG\[1\]
+ J2END_GH_BEG\[1\] J_l_GH_BEG\[1\] ConfigBits\[127\] ConfigBits\[128\] VGND VGND
+ VPWR VPWR B_ADR1 sky130_fd_sc_hd__mux4_2
XFILLER_0_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_ConfigMem_Inst_frame7_bit26 net67 net98 VGND VGND VPWR VPWR ConfigBits\[184\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1 AD0 AD1
+ AD2 AD3 ConfigBits\[110\] ConfigBits\[111\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XNN4END_inbuf_1__0_ net148 VGND VGND VPWR VPWR NN4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame7_bit15 net55 net98 VGND VGND VPWR VPWR ConfigBits\[173\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0951_ Inst_RegFile_32x4__1442_/Q Inst_RegFile_32x4__1438_/Q Inst_RegFile_32x4/_0335_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_cus_mux41_buf_inst1 J2END_CD_BEG\[3\]
+ JN2BEG\[5\] JS2BEG\[5\] JW2BEG\[5\] ConfigBits\[122\] ConfigBits\[123\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_A_ADR4_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1 net21
+ net161 net173 net214 ConfigBits\[330\] ConfigBits\[331\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0882_ Inst_RegFile_32x4/_0309_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0340_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1434_ net205 Inst_RegFile_32x4/_0086_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1434_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1296_ Inst_RegFile_32x4__1456_/Q Inst_RegFile_32x4/_0450_ Inst_RegFile_32x4/_0637_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0638_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1365_ net205 Inst_RegFile_32x4/_0025_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1365_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput486 net486 VGND VGND VPWR VPWR W6BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput453 net453 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput442 net442 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput431 net431 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput420 net420 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput464 net464 VGND VGND VPWR VPWR W2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput475 net475 VGND VGND VPWR VPWR W2BEGb[4] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_switch_matrix__04_ JE2BEG\[4\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__buf_1
Xoutput497 net497 VGND VGND VPWR VPWR WW4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_28__0_ FrameData_O_i\[28\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG1 net116 net16 net168
+ net221 ConfigBits\[192\] ConfigBits\[193\] VGND VGND VPWR VPWR J2MID_ABb_BEG\[1\]
+ sky130_fd_sc_hd__mux4_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[254\] ConfigBits\[255\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame3_bit21 net62 net94 VGND VGND VPWR VPWR ConfigBits\[307\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit10 net50 net94 VGND VGND VPWR VPWR ConfigBits\[296\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_D3 J2MID_ABa_BEG\[3\] J2MID_ABb_BEG\[3\]
+ J2END_AB_BEG\[3\] J_l_AB_BEG\[3\] ConfigBits\[142\] ConfigBits\[143\] VGND VGND
+ VPWR VPWR D3 sky130_fd_sc_hd__mux4_2
Xdata_outbuf_19__0_ FrameData_O_i\[19\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1150_ Inst_RegFile_32x4__1397_/Q Inst_RegFile_32x4/_0528_ Inst_RegFile_32x4/_0549_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1081_ Inst_RegFile_32x4__1361_/Q Inst_RegFile_32x4/_0496_ Inst_RegFile_32x4/_0508_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0510_ sky130_fd_sc_hd__mux2_1
XS4BEG_outbuf_8__0_ S4BEG_i\[8\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__0934_ Inst_RegFile_32x4__1406_/Q Inst_RegFile_32x4__1382_/Q Inst_RegFile_32x4/_0298_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0388_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0865_ Inst_RegFile_32x4__1344_/Q Inst_RegFile_32x4__1392_/Q Inst_RegFile_32x4__1464_/Q
+ Inst_RegFile_32x4__1460_/Q Inst_RegFile_32x4/_0321_ Inst_RegFile_32x4/_0322_ VGND
+ VGND VPWR VPWR Inst_RegFile_32x4/_0323_ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0796_ Inst_RegFile_32x4/_0173_ Inst_RegFile_32x4/_0258_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0259_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1279_ Inst_RegFile_32x4/_0628_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0100_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput283 net283 VGND VGND VPWR VPWR E6BEG[7] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1417_ net205 Inst_RegFile_32x4/_0069_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1417_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput294 net294 VGND VGND VPWR VPWR EE4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput272 net272 VGND VGND VPWR VPWR E2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput261 net261 VGND VGND VPWR VPWR E2BEG[3] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1348_ net205 Inst_RegFile_32x4/_0008_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1348_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame7_bit1 net60 net98 VGND VGND VPWR VPWR ConfigBits\[159\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2 net229
+ AD0 AD1 AD3 ConfigBits\[294\] ConfigBits\[295\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame6_bit25 net66 net97 VGND VGND VPWR VPWR ConfigBits\[215\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit14 net54 net97 VGND VGND VPWR VPWR ConfigBits\[204\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XS4END_inbuf_6__0_ net174 VGND VGND VPWR VPWR S4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1202_ Inst_RegFile_32x4/_0464_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0582_
+ sky130_fd_sc_hd__dlymetal6s2s_1
XInst_RegFile_32x4__1133_ Inst_RegFile_32x4/_0541_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0041_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1064_ Inst_RegFile_32x4/_0499_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0014_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0917_ Inst_RegFile_32x4__1441_/Q Inst_RegFile_32x4__1437_/Q Inst_RegFile_32x4/_0335_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0373_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0848_ Inst_RegFile_32x4/_0295_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0306_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame2_bit20 net61 net93 VGND VGND VPWR VPWR ConfigBits\[338\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0779_ Inst_RegFile_32x4/_0129_ Inst_RegFile_32x4/_0242_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0243_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_ConfigMem_Inst_frame2_bit31 net73 net93 VGND VGND VPWR VPWR ConfigBits\[349\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XEE4BEG_outbuf_7__0_ EE4BEG_i\[7\] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame9_bit18 net58 net100 VGND VGND VPWR VPWR ConfigBits\[112\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame9_bit29 net70 net100 VGND VGND VPWR VPWR ConfigBits\[123\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0702_ Inst_RegFile_32x4/_0134_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0168_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame5_bit24 net65 net96 VGND VGND VPWR VPWR ConfigBits\[246\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1116_ Inst_RegFile_32x4/_0531_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0034_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame5_bit13 net53 net96 VGND VGND VPWR VPWR ConfigBits\[235\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1047_ Inst_RegFile_32x4__1349_/Q Inst_RegFile_32x4/_0477_ Inst_RegFile_32x4/_0486_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0488_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame4_bit4 net75 net95 VGND VGND VPWR VPWR ConfigBits\[258\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst1 BD0 J2MID_EFa_BEG\[2\]
+ J2MID_GHa_BEG\[2\] J2END_AB_BEG\[2\] ConfigBits\[103\] ConfigBits\[104\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 J2MID_GHb_BEG\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2 net247
+ AD0 AD1 AD2 ConfigBits\[366\] ConfigBits\[367\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__1_/A1 ConfigBits\[96\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame1_bit30 net72 net92 VGND VGND VPWR VPWR ConfigBits\[380\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame8_bit28 net69 net99 VGND VGND VPWR VPWR ConfigBits\[154\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame8_bit17 net57 net99 VGND VGND VPWR VPWR ConfigBits\[143\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_S4BEG0 net24 net159 net180 AD0 ConfigBits\[66\]
+ ConfigBits\[67\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__mux4_1
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XNN4BEG_outbuf_11__0_ NN4BEG_i\[11\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_1
Xinput194 SS4END[14] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
Xinput183 S4END[4] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
Xinput172 S2MID[7] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_2
Xinput161 S2END[4] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_2
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput150 NN4END[7] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame4_bit23 net64 net95 VGND VGND VPWR VPWR ConfigBits\[277\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1 net12
+ net156 net164 net207 ConfigBits\[278\] ConfigBits\[279\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame4_bit12 net52 net95 VGND VGND VPWR VPWR ConfigBits\[266\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1450_ net205 Inst_RegFile_32x4/_0102_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1450_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1381_ net205 Inst_RegFile_32x4/_0041_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1381_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix__20_ JN2BEG\[4\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XNN4END_inbuf_10__0_ net142 VGND VGND VPWR VPWR NN4BEG_i\[10\] sky130_fd_sc_hd__buf_2
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_S1BEG3 BD3 J2MID_ABb_BEG\[2\] JE2BEG\[2\]
+ J_l_AB_BEG\[0\] ConfigBits\[64\] ConfigBits\[65\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__mux4_1
XFILLER_0_76_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame1_bit7 net78 net92 VGND VGND VPWR VPWR ConfigBits\[357\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_ConfigMem_Inst_frame11_bit3 net74 net83 VGND VGND VPWR VPWR ConfigBits\[33\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR W_ADR4 sky130_fd_sc_hd__buf_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst1 BD2 J2MID_ABa_BEG\[2\]
+ J2MID_CDa_BEG\[2\] J2END_EF_BEG\[3\] ConfigBits\[77\] ConfigBits\[78\] VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__1_/A1
+ sky130_fd_sc_hd__mux4_1
Xstrobe_outbuf_11__0_ FrameStrobe_O_i\[11\] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_6__0_ FrameData_O_i\[6\] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_B_ADR2 J2MID_GHa_BEG\[2\] J2MID_GHb_BEG\[2\]
+ J2END_GH_BEG\[2\] J_l_GH_BEG\[2\] ConfigBits\[129\] ConfigBits\[130\] VGND VGND
+ VPWR VPWR B_ADR2 sky130_fd_sc_hd__mux4_2
XFILLER_0_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame7_bit16 net56 net98 VGND VGND VPWR VPWR ConfigBits\[174\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame7_bit27 net68 net98 VGND VGND VPWR VPWR ConfigBits\[185\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2 BD0 BD1
+ BD2 BD3 ConfigBits\[110\] ConfigBits\[111\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_32x4__0950_ Inst_RegFile_32x4/_0329_ Inst_RegFile_32x4/_0403_ Inst_RegFile_32x4/_0319_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0404_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0881_ Inst_RegFile_32x4__1432_/Q Inst_RegFile_32x4__1428_/Q Inst_RegFile_32x4/_0338_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0339_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2 net226
+ AD0 AD1 AD2 ConfigBits\[330\] ConfigBits\[331\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__1433_ net205 Inst_RegFile_32x4/_0085_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1433_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1295_ Inst_RegFile_32x4/_0473_ Inst_RegFile_32x4/_0626_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0637_ sky130_fd_sc_hd__nor2_2
XInst_RegFile_switch_matrix__03_ JE2BEG\[3\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__buf_1
XInst_RegFile_32x4__1364_ net205 Inst_RegFile_32x4/_0024_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1364_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput487 net487 VGND VGND VPWR VPWR W6BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput443 net443 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput454 net454 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput432 net432 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput410 net410 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput421 net421 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput465 net465 VGND VGND VPWR VPWR W2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput476 net476 VGND VGND VPWR VPWR W2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput498 net498 VGND VGND VPWR VPWR WW4BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XWW4END_inbuf_2__0_ net250 VGND VGND VPWR VPWR WW4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG2 net118 net18 net170
+ net223 ConfigBits\[194\] ConfigBits\[195\] VGND VGND VPWR VPWR J2MID_ABb_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_20_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xstrobe_inbuf_9__0_ net100 VGND VGND VPWR VPWR FrameStrobe_O_i\[9\] sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3/X ConfigBits\[256\]
+ ConfigBits\[257\] VGND VGND VPWR VPWR JN2BEG\[0\] sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame3_bit22 net63 net94 VGND VGND VPWR VPWR ConfigBits\[308\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit11 net51 net94 VGND VGND VPWR VPWR ConfigBits\[297\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1080_ Inst_RegFile_32x4/_0509_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0020_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0933_ Inst_RegFile_32x4/_0290_ Inst_RegFile_32x4/_0386_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0387_ sky130_fd_sc_hd__and2b_1
XInst_RegFile_32x4__0864_ B_ADR1 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0322_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1416_ net205 Inst_RegFile_32x4/_0068_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1416_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__0795_ Inst_RegFile_32x4__1379_/Q Inst_RegFile_32x4__1375_/Q Inst_RegFile_32x4/_0174_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1278_ Inst_RegFile_32x4__1448_/Q Inst_RegFile_32x4/_0591_ Inst_RegFile_32x4/_0627_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0628_ sky130_fd_sc_hd__mux2_1
Xoutput284 net284 VGND VGND VPWR VPWR E6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput295 net295 VGND VGND VPWR VPWR EE4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput273 net273 VGND VGND VPWR VPWR E2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput262 net262 VGND VGND VPWR VPWR E2BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__1347_ net205 Inst_RegFile_32x4/_0007_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1347_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[294\] ConfigBits\[295\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame7_bit2 net71 net98 VGND VGND VPWR VPWR ConfigBits\[160\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame6_bit26 net67 net97 VGND VGND VPWR VPWR ConfigBits\[216\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit15 net55 net97 VGND VGND VPWR VPWR ConfigBits\[205\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1201_ Inst_RegFile_32x4/_0581_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0069_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_32x4__1132_ Inst_RegFile_32x4__1381_/Q Inst_RegFile_32x4/_0528_ Inst_RegFile_32x4/_0539_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0541_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1063_ Inst_RegFile_32x4__1354_/Q Inst_RegFile_32x4/_0498_ Inst_RegFile_32x4/_0494_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0778_ Inst_RegFile_32x4__1442_/Q Inst_RegFile_32x4__1438_/Q Inst_RegFile_32x4/_0174_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0242_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0916_ Inst_RegFile_32x4/_0329_ Inst_RegFile_32x4/_0371_ Inst_RegFile_32x4/_0332_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0372_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0847_ Inst_RegFile_32x4/_0302_ Inst_RegFile_32x4/_0304_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0305_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame2_bit21 net62 net93 VGND VGND VPWR VPWR ConfigBits\[339\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame2_bit10 net50 net93 VGND VGND VPWR VPWR ConfigBits\[328\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame9_bit19 net59 net100 VGND VGND VPWR VPWR ConfigBits\[113\]
+ Inst_RegFile_ConfigMem_Inst_frame9_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XE6END_inbuf_2__0_ net27 VGND VGND VPWR VPWR E6BEG_i\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_32x4__0701_ Inst_RegFile_32x4/_0152_ Inst_RegFile_32x4/_0166_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0167_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame5_bit25 net66 net96 VGND VGND VPWR VPWR ConfigBits\[247\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1115_ Inst_RegFile_32x4__1374_/Q Inst_RegFile_32x4/_0530_ Inst_RegFile_32x4/_0526_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0531_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame5_bit14 net54 net96 VGND VGND VPWR VPWR ConfigBits\[236\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1046_ Inst_RegFile_32x4/_0487_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0008_
+ sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame4_bit5 net76 net95 VGND VGND VPWR VPWR ConfigBits\[259\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XSS4END_inbuf_4__0_ net203 VGND VGND VPWR VPWR SS4BEG_i\[4\] sky130_fd_sc_hd__buf_2
XFILLER_0_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_3 J2MID_GHb_BEG\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3 AD3 BD1
+ BD2 BD3 ConfigBits\[366\] ConfigBits\[367\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_6__0_ FrameStrobe_O_i\[6\] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame1_bit20 net61 net92 VGND VGND VPWR VPWR ConfigBits\[370\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame1_bit31 net73 net92 VGND VGND VPWR VPWR ConfigBits\[381\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame8_bit18 net58 net99 VGND VGND VPWR VPWR ConfigBits\[144\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame8_bit29 net70 net99 VGND VGND VPWR VPWR ConfigBits\[155\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_S4BEG1 net21 net160 net181 AD1 ConfigBits\[68\]
+ ConfigBits\[69\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__mux4_1
XInst_RegFile_32x4__1029_ Inst_RegFile_32x4/_0471_ Inst_RegFile_32x4/_0474_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0475_ sky130_fd_sc_hd__and2_2
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XEE4END_inbuf_3__0_ net46 VGND VGND VPWR VPWR EE4BEG_i\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_0__0_ net49 VGND VGND VPWR VPWR FrameData_O_i\[0\] sky130_fd_sc_hd__buf_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput162 S2END[5] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_2
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput151 NN4END[8] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
Xinput140 NN4END[12] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
Xinput195 SS4END[15] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
Xinput184 S4END[5] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xinput173 S4END[0] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_4
XWW4BEG_outbuf_4__0_ WW4BEG_i\[4\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2 net209
+ AD0 AD1 AD2 ConfigBits\[278\] ConfigBits\[279\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame4_bit24 net65 net95 VGND VGND VPWR VPWR ConfigBits\[278\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_ConfigMem_Inst_frame4_bit13 net53 net95 VGND VGND VPWR VPWR ConfigBits\[267\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1380_ net205 Inst_RegFile_32x4/_0040_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1380_/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_ConfigMem_Inst_frame1_bit8 net79 net92 VGND VGND VPWR VPWR ConfigBits\[358\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_my_mux2_inst__1_/A1 ConfigBits\[154\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_W_ADR4_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XInst_RegFile_ConfigMem_Inst_frame11_bit4 net75 net83 VGND VGND VPWR VPWR ConfigBits\[34\]
+ Inst_RegFile_ConfigMem_Inst_frame11_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XE6BEG_outbuf_7__0_ E6BEG_i\[7\] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_B_ADR3 J2MID_GHa_BEG\[3\] J2MID_GHb_BEG\[3\]
+ J2END_GH_BEG\[3\] J_l_GH_BEG\[3\] ConfigBits\[131\] ConfigBits\[132\] VGND VGND
+ VPWR VPWR B_ADR3 sky130_fd_sc_hd__mux4_2
XInst_RegFile_ConfigMem_Inst_frame0_bit30 net72 net81 VGND VGND VPWR VPWR ConfigBits\[412\]
+ Inst_RegFile_ConfigMem_Inst_frame0_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame7_bit17 net57 net98 VGND VGND VPWR VPWR ConfigBits\[175\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3 J2MID_ABa_BEG\[2\]
+ J2MID_CDa_BEG\[2\] J2MID_EFa_BEG\[2\] J2MID_GHa_BEG\[2\] ConfigBits\[110\] ConfigBits\[111\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame7_bit28 net69 net98 VGND VGND VPWR VPWR ConfigBits\[186\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3 BD0 BD1
+ BD2 BD3 ConfigBits\[330\] ConfigBits\[331\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_32x4__0880_ Inst_RegFile_32x4/_0297_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0338_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput400 net400 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1432_ net205 Inst_RegFile_32x4/_0084_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1432_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput411 net411 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__clkbuf_4
XN4END_inbuf_6__0_ net122 VGND VGND VPWR VPWR N4BEG_i\[6\] sky130_fd_sc_hd__buf_2
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1294_ Inst_RegFile_32x4/_0636_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0107_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_switch_matrix__02_ JE2BEG\[2\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_1
Xoutput488 net488 VGND VGND VPWR VPWR W6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput444 net444 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput455 net455 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput433 net433 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput422 net422 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput466 net466 VGND VGND VPWR VPWR W2BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1363_ net205 Inst_RegFile_32x4/_0023_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1363_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput477 net477 VGND VGND VPWR VPWR W2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput499 net499 VGND VGND VPWR VPWR WW4BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG3 net114 net14 net166
+ net219 ConfigBits\[196\] ConfigBits\[197\] VGND VGND VPWR VPWR J2MID_ABb_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame3_bit23 net64 net94 VGND VGND VPWR VPWR ConfigBits\[309\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame3_bit12 net52 net94 VGND VGND VPWR VPWR ConfigBits\[298\]
+ Inst_RegFile_ConfigMem_Inst_frame3_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0932_ Inst_RegFile_32x4__1358_/Q Inst_RegFile_32x4__1446_/Q Inst_RegFile_32x4/_0292_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0386_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__0794_ Inst_RegFile_32x4/_0185_ Inst_RegFile_32x4/_0256_ Inst_RegFile_32x4/_0139_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0257_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_32x4__0863_ Inst_RegFile_32x4/_0297_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0321_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__1415_ net205 Inst_RegFile_32x4/_0067_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1415_/Q
+ sky130_fd_sc_hd__dfxtp_1
XInst_RegFile_32x4__1346_ net205 Inst_RegFile_32x4/_0006_ VGND VGND VPWR VPWR Inst_RegFile_32x4__1346_/Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput285 net285 VGND VGND VPWR VPWR E6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput274 net274 VGND VGND VPWR VPWR E6BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput296 net296 VGND VGND VPWR VPWR EE4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput263 net263 VGND VGND VPWR VPWR E2BEG[5] sky130_fd_sc_hd__clkbuf_4
XInst_RegFile_32x4__1277_ Inst_RegFile_32x4/_0493_ Inst_RegFile_32x4/_0626_ VGND VGND
+ VPWR VPWR Inst_RegFile_32x4/_0627_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3/X ConfigBits\[296\]
+ ConfigBits\[297\] VGND VGND VPWR VPWR JE2BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame7_bit3 net74 net98 VGND VGND VPWR VPWR ConfigBits\[161\]
+ Inst_RegFile_ConfigMem_Inst_frame7_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame6_bit16 net56 net97 VGND VGND VPWR VPWR ConfigBits\[206\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_33_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_ConfigMem_Inst_frame6_bit27 net68 net97 VGND VGND VPWR VPWR ConfigBits\[217\]
+ Inst_RegFile_ConfigMem_Inst_frame6_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1200_ Inst_RegFile_32x4/_0580_ Inst_RegFile_32x4__1417_/Q Inst_RegFile_32x4/_0578_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__1_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__1_/A0
+ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__1_/A1 ConfigBits\[85\]
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1062_ Inst_RegFile_32x4/_0464_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0498_
+ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_32x4__1131_ Inst_RegFile_32x4/_0540_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0040_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RegFile_32x4__0915_ Inst_RegFile_32x4__1449_/Q Inst_RegFile_32x4__1473_/Q Inst_RegFile_32x4/_0317_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_ConfigMem_Inst_frame2_bit22 net63 net93 VGND VGND VPWR VPWR ConfigBits\[340\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RegFile_32x4__0777_ Inst_RegFile_32x4/_0168_ Inst_RegFile_32x4/_0240_ Inst_RegFile_32x4/_0158_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0241_ sky130_fd_sc_hd__a21o_1
XInst_RegFile_ConfigMem_Inst_frame2_bit11 net51 net93 VGND VGND VPWR VPWR ConfigBits\[329\]
+ Inst_RegFile_ConfigMem_Inst_frame2_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__0846_ Inst_RegFile_32x4__1376_/Q Inst_RegFile_32x4__1372_/Q Inst_RegFile_32x4/_0303_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__1329_ Inst_RegFile_32x4/_0481_ Inst_RegFile_32x4__1471_/Q Inst_RegFile_32x4/_0652_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_my_mux2_inst__2_ Inst_RegFile_switch_matrix_inst_cus_mux81_buf_B_ADR4_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR B_ADR4 sky130_fd_sc_hd__buf_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_32x4__0700_ Inst_RegFile_32x4__1456_/Q Inst_RegFile_32x4__1452_/Q Inst_RegFile_32x4/_0165_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0166_ sky130_fd_sc_hd__mux2_1
XNN4BEG_outbuf_7__0_ NN4BEG_i\[7\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_1
XInst_RegFile_ConfigMem_Inst_frame5_bit26 net67 net96 VGND VGND VPWR VPWR ConfigBits\[248\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame5_bit15 net55 net96 VGND VGND VPWR VPWR ConfigBits\[237\]
+ Inst_RegFile_ConfigMem_Inst_frame5_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_32x4__1045_ Inst_RegFile_32x4__1348_/Q Inst_RegFile_32x4/_0470_ Inst_RegFile_32x4/_0486_
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0487_ sky130_fd_sc_hd__mux2_1
XInst_RegFile_32x4__1114_ D2 VGND VGND VPWR VPWR Inst_RegFile_32x4/_0530_ sky130_fd_sc_hd__clkbuf_2
XInst_RegFile_ConfigMem_Inst_frame4_bit6 net77 net95 VGND VGND VPWR VPWR ConfigBits\[260\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RegFile_32x4__0829_ Inst_RegFile_32x4__1387_/D Inst_RegFile_32x4__1387_/Q ConfigBits\[0\]
+ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 JN2BEG\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst4 Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1/X Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2/X
+ Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3/X ConfigBits\[368\]
+ ConfigBits\[369\] VGND VGND VPWR VPWR JW2BEG\[4\] sky130_fd_sc_hd__mux4_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RegFile_ConfigMem_Inst_frame1_bit21 net62 net92 VGND VGND VPWR VPWR ConfigBits\[371\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame8_bit19 net59 net99 VGND VGND VPWR VPWR ConfigBits\[145\]
+ Inst_RegFile_ConfigMem_Inst_frame8_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RegFile_ConfigMem_Inst_frame1_bit10 net50 net92 VGND VGND VPWR VPWR ConfigBits\[360\]
+ Inst_RegFile_ConfigMem_Inst_frame1_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RegFile_switch_matrix_inst_cus_mux41_buf_S4BEG2 net157 net182 net229 AD2 ConfigBits\[70\]
+ ConfigBits\[71\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__mux4_2
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_32x4__1028_ Inst_RegFile_32x4/_0473_ VGND VGND VPWR VPWR Inst_RegFile_32x4/_0474_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput196 SS4END[1] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_4
Xinput174 S4END[10] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
Xinput185 S4END[6] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
Xinput163 S2END[6] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xinput141 NN4END[13] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
Xinput152 NN4END[9] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
Xinput130 N4END[3] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_2
XFILLER_0_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3 AD3 BD0
+ BD1 BD3 ConfigBits\[278\] ConfigBits\[279\] VGND VGND VPWR VPWR Inst_RegFile_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_RegFile_ConfigMem_Inst_frame4_bit25 net66 net95 VGND VGND VPWR VPWR ConfigBits\[279\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RegFile_ConfigMem_Inst_frame4_bit14 net54 net95 VGND VGND VPWR VPWR ConfigBits\[268\]
+ Inst_RegFile_ConfigMem_Inst_frame4_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XNN4END_inbuf_4__0_ net151 VGND VGND VPWR VPWR NN4BEG_i\[4\] sky130_fd_sc_hd__clkbuf_2
.ends

