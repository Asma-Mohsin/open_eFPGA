magic
tech sky130A
magscale 1 2
timestamp 1733306926
<< viali >>
rect 1777 8585 1811 8619
rect 2697 8585 2731 8619
rect 3065 8585 3099 8619
rect 3433 8585 3467 8619
rect 3985 8585 4019 8619
rect 4537 8585 4571 8619
rect 5089 8585 5123 8619
rect 5641 8585 5675 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7113 8585 7147 8619
rect 8033 8585 8067 8619
rect 8585 8585 8619 8619
rect 9045 8585 9079 8619
rect 10057 8585 10091 8619
rect 10609 8585 10643 8619
rect 11161 8585 11195 8619
rect 11713 8585 11747 8619
rect 12265 8585 12299 8619
rect 12817 8585 12851 8619
rect 13737 8585 13771 8619
rect 14657 8585 14691 8619
rect 15025 8585 15059 8619
rect 15761 8585 15795 8619
rect 16313 8585 16347 8619
rect 17049 8585 17083 8619
rect 17601 8585 17635 8619
rect 18061 8585 18095 8619
rect 18613 8585 18647 8619
rect 18981 8585 19015 8619
rect 20177 8585 20211 8619
rect 22937 8585 22971 8619
rect 24041 8585 24075 8619
rect 30665 8585 30699 8619
rect 31769 8585 31803 8619
rect 32137 8585 32171 8619
rect 32505 8585 32539 8619
rect 33241 8585 33275 8619
rect 33609 8585 33643 8619
rect 33977 8585 34011 8619
rect 34713 8585 34747 8619
rect 35449 8585 35483 8619
rect 36185 8585 36219 8619
rect 36553 8585 36587 8619
rect 38025 8585 38059 8619
rect 39129 8585 39163 8619
rect 40049 8585 40083 8619
rect 40601 8585 40635 8619
rect 41521 8585 41555 8619
rect 42625 8585 42659 8619
rect 44281 8585 44315 8619
rect 45753 8585 45787 8619
rect 2789 8517 2823 8551
rect 5181 8517 5215 8551
rect 5733 8517 5767 8551
rect 9413 8517 9447 8551
rect 9781 8517 9815 8551
rect 10701 8517 10735 8551
rect 19257 8517 19291 8551
rect 43085 8517 43119 8551
rect 45661 8517 45695 8551
rect 1961 8449 1995 8483
rect 2329 8449 2363 8483
rect 3249 8449 3283 8483
rect 3617 8449 3651 8483
rect 4261 8449 4295 8483
rect 4721 8449 4755 8483
rect 6193 8449 6227 8483
rect 6837 8449 6871 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 8125 8449 8159 8483
rect 8677 8449 8711 8483
rect 9229 8449 9263 8483
rect 10241 8449 10275 8483
rect 11253 8449 11287 8483
rect 11897 8449 11931 8483
rect 12357 8449 12391 8483
rect 13001 8449 13035 8483
rect 13369 8449 13403 8483
rect 13829 8449 13863 8483
rect 14749 8449 14783 8483
rect 15301 8449 15335 8483
rect 15957 8449 15991 8483
rect 16405 8449 16439 8483
rect 17233 8449 17267 8483
rect 17693 8449 17727 8483
rect 17969 8449 18003 8483
rect 18429 8449 18463 8483
rect 18797 8449 18831 8483
rect 19625 8449 19659 8483
rect 19993 8449 20027 8483
rect 20361 8449 20395 8483
rect 21097 8449 21131 8483
rect 21373 8449 21407 8483
rect 21649 8449 21683 8483
rect 22017 8449 22051 8483
rect 22293 8449 22327 8483
rect 22385 8449 22419 8483
rect 22845 8449 22879 8483
rect 23121 8449 23155 8483
rect 23397 8449 23431 8483
rect 23673 8449 23707 8483
rect 23949 8449 23983 8483
rect 24225 8449 24259 8483
rect 24593 8449 24627 8483
rect 24961 8449 24995 8483
rect 25329 8449 25363 8483
rect 25697 8449 25731 8483
rect 26065 8449 26099 8483
rect 26433 8449 26467 8483
rect 26801 8449 26835 8483
rect 27169 8449 27203 8483
rect 27537 8449 27571 8483
rect 27905 8449 27939 8483
rect 28273 8449 28307 8483
rect 28641 8449 28675 8483
rect 29009 8449 29043 8483
rect 29377 8449 29411 8483
rect 29745 8449 29779 8483
rect 30113 8449 30147 8483
rect 30481 8449 30515 8483
rect 30849 8449 30883 8483
rect 31217 8449 31251 8483
rect 31585 8449 31619 8483
rect 31953 8449 31987 8483
rect 32321 8449 32355 8483
rect 32689 8449 32723 8483
rect 33057 8449 33091 8483
rect 33425 8449 33459 8483
rect 33793 8449 33827 8483
rect 34161 8449 34195 8483
rect 34529 8449 34563 8483
rect 34897 8449 34931 8483
rect 35265 8449 35299 8483
rect 35633 8449 35667 8483
rect 36001 8449 36035 8483
rect 36369 8449 36403 8483
rect 36737 8449 36771 8483
rect 37105 8449 37139 8483
rect 37473 8449 37507 8483
rect 37841 8449 37875 8483
rect 38209 8449 38243 8483
rect 38577 8449 38611 8483
rect 38945 8449 38979 8483
rect 39313 8449 39347 8483
rect 39957 8449 39991 8483
rect 40509 8449 40543 8483
rect 40969 8449 41003 8483
rect 41429 8449 41463 8483
rect 42533 8449 42567 8483
rect 43637 8449 43671 8483
rect 44189 8449 44223 8483
rect 45109 8449 45143 8483
rect 45385 8381 45419 8415
rect 2145 8313 2179 8347
rect 7481 8313 7515 8347
rect 13185 8313 13219 8347
rect 20545 8313 20579 8347
rect 23489 8313 23523 8347
rect 24409 8313 24443 8347
rect 26249 8313 26283 8347
rect 27721 8313 27755 8347
rect 28089 8313 28123 8347
rect 32873 8313 32907 8347
rect 34345 8313 34379 8347
rect 35081 8313 35115 8347
rect 35817 8313 35851 8347
rect 36921 8313 36955 8347
rect 38393 8313 38427 8347
rect 38761 8313 38795 8347
rect 41153 8313 41187 8347
rect 43269 8313 43303 8347
rect 43821 8313 43855 8347
rect 20913 8245 20947 8279
rect 21189 8245 21223 8279
rect 21465 8245 21499 8279
rect 21833 8245 21867 8279
rect 22109 8245 22143 8279
rect 22569 8245 22603 8279
rect 22661 8245 22695 8279
rect 23213 8245 23247 8279
rect 23765 8245 23799 8279
rect 24777 8245 24811 8279
rect 25145 8245 25179 8279
rect 25513 8245 25547 8279
rect 25881 8245 25915 8279
rect 26617 8245 26651 8279
rect 26985 8245 27019 8279
rect 27353 8245 27387 8279
rect 28457 8245 28491 8279
rect 28825 8245 28859 8279
rect 29193 8245 29227 8279
rect 29561 8245 29595 8279
rect 29929 8245 29963 8279
rect 30297 8245 30331 8279
rect 31033 8245 31067 8279
rect 31401 8245 31435 8279
rect 37289 8245 37323 8279
rect 37657 8245 37691 8279
rect 1869 8041 1903 8075
rect 4077 8041 4111 8075
rect 4629 8041 4663 8075
rect 6653 8041 6687 8075
rect 7205 8041 7239 8075
rect 9229 8041 9263 8075
rect 10057 8041 10091 8075
rect 11805 8041 11839 8075
rect 12633 8041 12667 8075
rect 14381 8041 14415 8075
rect 14933 8041 14967 8075
rect 15577 8041 15611 8075
rect 17049 8041 17083 8075
rect 17785 8041 17819 8075
rect 18061 8041 18095 8075
rect 18337 8041 18371 8075
rect 18797 8041 18831 8075
rect 19625 8041 19659 8075
rect 19901 8041 19935 8075
rect 20453 8041 20487 8075
rect 20729 8041 20763 8075
rect 21005 8041 21039 8075
rect 21281 8041 21315 8075
rect 21833 8041 21867 8075
rect 23765 8041 23799 8075
rect 24501 8041 24535 8075
rect 25421 8041 25455 8075
rect 25697 8041 25731 8075
rect 27721 8041 27755 8075
rect 28089 8041 28123 8075
rect 28457 8041 28491 8075
rect 29653 8041 29687 8075
rect 41153 8041 41187 8075
rect 43361 8041 43395 8075
rect 45201 8041 45235 8075
rect 45937 8041 45971 8075
rect 2421 7973 2455 8007
rect 22661 7973 22695 8007
rect 24041 7973 24075 8007
rect 26525 7973 26559 8007
rect 27077 7973 27111 8007
rect 44189 7973 44223 8007
rect 2605 7837 2639 7871
rect 4813 7837 4847 7871
rect 7389 7837 7423 7871
rect 10241 7837 10275 7871
rect 12817 7837 12851 7871
rect 15117 7837 15151 7871
rect 15761 7837 15795 7871
rect 17233 7837 17267 7871
rect 17969 7837 18003 7871
rect 18245 7837 18279 7871
rect 18521 7837 18555 7871
rect 18613 7837 18647 7871
rect 19073 7837 19107 7871
rect 19533 7837 19567 7871
rect 19809 7837 19843 7871
rect 20085 7837 20119 7871
rect 20361 7837 20395 7871
rect 20637 7837 20671 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 21465 7837 21499 7871
rect 21741 7837 21775 7871
rect 22017 7837 22051 7871
rect 22293 7837 22327 7871
rect 22569 7837 22603 7871
rect 22845 7837 22879 7871
rect 23121 7837 23155 7871
rect 23397 7837 23431 7871
rect 23673 7837 23707 7871
rect 23949 7837 23983 7871
rect 24225 7837 24259 7871
rect 24685 7837 24719 7871
rect 24961 7837 24995 7871
rect 25329 7837 25363 7871
rect 25605 7837 25639 7871
rect 25881 7837 25915 7871
rect 26157 7837 26191 7871
rect 26433 7837 26467 7871
rect 26709 7837 26743 7871
rect 26985 7837 27019 7871
rect 27261 7837 27295 7871
rect 27537 7837 27571 7871
rect 27905 7837 27939 7871
rect 28273 7837 28307 7871
rect 28641 7837 28675 7871
rect 29009 7837 29043 7871
rect 29377 7837 29411 7871
rect 29837 7837 29871 7871
rect 40969 7837 41003 7871
rect 2145 7769 2179 7803
rect 4353 7769 4387 7803
rect 6929 7769 6963 7803
rect 9505 7769 9539 7803
rect 12081 7769 12115 7803
rect 14657 7769 14691 7803
rect 43269 7769 43303 7803
rect 44005 7769 44039 7803
rect 45109 7769 45143 7803
rect 45661 7769 45695 7803
rect 18889 7701 18923 7735
rect 19349 7701 19383 7735
rect 20177 7701 20211 7735
rect 21557 7701 21591 7735
rect 22109 7701 22143 7735
rect 22385 7701 22419 7735
rect 22937 7701 22971 7735
rect 23213 7701 23247 7735
rect 23489 7701 23523 7735
rect 24777 7701 24811 7735
rect 25145 7701 25179 7735
rect 25973 7701 26007 7735
rect 26249 7701 26283 7735
rect 26801 7701 26835 7735
rect 27353 7701 27387 7735
rect 28825 7701 28859 7735
rect 29193 7701 29227 7735
rect 1501 7497 1535 7531
rect 20177 7497 20211 7531
rect 20637 7497 20671 7531
rect 22569 7497 22603 7531
rect 23121 7497 23155 7531
rect 24685 7497 24719 7531
rect 45109 7497 45143 7531
rect 45661 7497 45695 7531
rect 46397 7497 46431 7531
rect 44833 7429 44867 7463
rect 1777 7361 1811 7395
rect 19809 7361 19843 7395
rect 19993 7361 20027 7395
rect 20545 7361 20579 7395
rect 20821 7361 20855 7395
rect 22753 7361 22787 7395
rect 23305 7361 23339 7395
rect 23581 7361 23615 7395
rect 23857 7361 23891 7395
rect 24225 7361 24259 7395
rect 24593 7361 24627 7395
rect 24869 7361 24903 7395
rect 44465 7361 44499 7395
rect 45017 7361 45051 7395
rect 45569 7361 45603 7395
rect 46121 7361 46155 7395
rect 23673 7225 23707 7259
rect 19625 7157 19659 7191
rect 20361 7157 20395 7191
rect 23397 7157 23431 7191
rect 24041 7157 24075 7191
rect 24409 7157 24443 7191
rect 46213 6953 46247 6987
rect 45845 6817 45879 6851
rect 46121 6749 46155 6783
rect 45569 6681 45603 6715
rect 23673 2601 23707 2635
rect 24225 2601 24259 2635
rect 24777 2601 24811 2635
rect 25605 2601 25639 2635
rect 27721 2601 27755 2635
rect 29929 2601 29963 2635
rect 32137 2601 32171 2635
rect 34345 2601 34379 2635
rect 38853 2601 38887 2635
rect 43269 2601 43303 2635
rect 45201 2601 45235 2635
rect 45661 2601 45695 2635
rect 45753 2601 45787 2635
rect 25053 2533 25087 2567
rect 25329 2533 25363 2567
rect 36645 2533 36679 2567
rect 23397 2465 23431 2499
rect 23489 2397 23523 2431
rect 23765 2397 23799 2431
rect 24041 2397 24075 2431
rect 24593 2397 24627 2431
rect 24869 2397 24903 2431
rect 25145 2397 25179 2431
rect 25421 2397 25455 2431
rect 27537 2397 27571 2431
rect 29745 2397 29779 2431
rect 31953 2397 31987 2431
rect 34161 2397 34195 2431
rect 36461 2397 36495 2431
rect 38669 2397 38703 2431
rect 43085 2397 43119 2431
rect 45017 2397 45051 2431
rect 45477 2397 45511 2431
rect 45937 2397 45971 2431
rect 21097 2329 21131 2363
rect 23213 2329 23247 2363
rect 21189 2261 21223 2295
rect 23949 2261 23983 2295
rect 20269 2057 20303 2091
rect 22385 2057 22419 2091
rect 22661 2057 22695 2091
rect 23397 2057 23431 2091
rect 23949 2057 23983 2091
rect 24685 2057 24719 2091
rect 27169 2057 27203 2091
rect 29285 2057 29319 2091
rect 31401 2057 31435 2091
rect 33701 2057 33735 2091
rect 35725 2057 35759 2091
rect 37933 2057 37967 2091
rect 42625 2057 42659 2091
rect 44281 2057 44315 2091
rect 45845 2057 45879 2091
rect 20085 1921 20119 1955
rect 22201 1921 22235 1955
rect 22477 1921 22511 1955
rect 22937 1921 22971 1955
rect 23213 1921 23247 1955
rect 23489 1921 23523 1955
rect 23765 1921 23799 1955
rect 24041 1921 24075 1955
rect 24501 1921 24535 1955
rect 24777 1921 24811 1955
rect 26985 1921 27019 1955
rect 29101 1921 29135 1955
rect 31217 1921 31251 1955
rect 33517 1921 33551 1955
rect 35541 1921 35575 1955
rect 37749 1921 37783 1955
rect 42441 1921 42475 1955
rect 44097 1921 44131 1955
rect 44557 1921 44591 1955
rect 45661 1921 45695 1955
rect 23121 1785 23155 1819
rect 44741 1785 44775 1819
rect 23673 1717 23707 1751
rect 24225 1717 24259 1751
rect 24961 1717 24995 1751
rect 19809 1513 19843 1547
rect 22017 1513 22051 1547
rect 23673 1513 23707 1547
rect 24225 1513 24259 1547
rect 26433 1513 26467 1547
rect 28641 1513 28675 1547
rect 30849 1513 30883 1547
rect 33057 1513 33091 1547
rect 35265 1513 35299 1547
rect 37473 1513 37507 1547
rect 41889 1513 41923 1547
rect 44097 1513 44131 1547
rect 46121 1513 46155 1547
rect 15393 1445 15427 1479
rect 23397 1445 23431 1479
rect 1961 1309 1995 1343
rect 4169 1309 4203 1343
rect 6377 1309 6411 1343
rect 8585 1309 8619 1343
rect 10793 1309 10827 1343
rect 13001 1309 13035 1343
rect 15209 1309 15243 1343
rect 17417 1309 17451 1343
rect 19625 1309 19659 1343
rect 21833 1309 21867 1343
rect 23213 1309 23247 1343
rect 23489 1309 23523 1343
rect 24041 1309 24075 1343
rect 26249 1309 26283 1343
rect 28457 1309 28491 1343
rect 30665 1309 30699 1343
rect 32873 1309 32907 1343
rect 35081 1309 35115 1343
rect 37289 1309 37323 1343
rect 39497 1309 39531 1343
rect 41705 1309 41739 1343
rect 43913 1309 43947 1343
rect 46305 1309 46339 1343
rect 2145 1173 2179 1207
rect 4353 1173 4387 1207
rect 6561 1173 6595 1207
rect 8769 1173 8803 1207
rect 10977 1173 11011 1207
rect 13185 1173 13219 1207
rect 17601 1173 17635 1207
rect 39681 1173 39715 1207
<< metal1 >>
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 16850 9976 16856 9988
rect 7248 9948 16856 9976
rect 7248 9936 7254 9948
rect 16850 9936 16856 9948
rect 16908 9936 16914 9988
rect 21542 9976 21548 9988
rect 17052 9948 21548 9976
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 17052 9908 17080 9948
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 24026 9936 24032 9988
rect 24084 9976 24090 9988
rect 35066 9976 35072 9988
rect 24084 9948 35072 9976
rect 24084 9936 24090 9948
rect 35066 9936 35072 9948
rect 35124 9936 35130 9988
rect 20714 9908 20720 9920
rect 10192 9880 17080 9908
rect 17144 9880 20720 9908
rect 10192 9868 10198 9880
rect 12710 9800 12716 9852
rect 12768 9840 12774 9852
rect 16114 9840 16120 9852
rect 12768 9812 16120 9840
rect 12768 9800 12774 9812
rect 16114 9800 16120 9812
rect 16172 9800 16178 9852
rect 17144 9772 17172 9880
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 20898 9868 20904 9920
rect 20956 9908 20962 9920
rect 22278 9908 22284 9920
rect 20956 9880 22284 9908
rect 20956 9868 20962 9880
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 28810 9908 28816 9920
rect 24320 9880 28816 9908
rect 22186 9840 22192 9852
rect 6196 9744 17172 9772
rect 17236 9812 22192 9840
rect 6196 9648 6224 9744
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 17236 9704 17264 9812
rect 22186 9800 22192 9812
rect 22244 9800 22250 9852
rect 24320 9840 24348 9880
rect 28810 9868 28816 9880
rect 28868 9868 28874 9920
rect 28902 9868 28908 9920
rect 28960 9908 28966 9920
rect 28960 9880 31754 9908
rect 28960 9868 28966 9880
rect 22480 9812 24348 9840
rect 17402 9732 17408 9784
rect 17460 9772 17466 9784
rect 22480 9772 22508 9812
rect 24394 9800 24400 9852
rect 24452 9840 24458 9852
rect 24452 9812 29408 9840
rect 24452 9800 24458 9812
rect 27062 9772 27068 9784
rect 17460 9744 22508 9772
rect 22572 9744 27068 9772
rect 17460 9732 17466 9744
rect 11940 9676 17264 9704
rect 11940 9664 11946 9676
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 22572 9704 22600 9744
rect 27062 9732 27068 9744
rect 27120 9732 27126 9784
rect 17920 9676 22600 9704
rect 17920 9664 17926 9676
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 24210 9704 24216 9716
rect 22704 9676 24216 9704
rect 22704 9664 22710 9676
rect 24210 9664 24216 9676
rect 24268 9664 24274 9716
rect 29270 9704 29276 9716
rect 28966 9676 29276 9704
rect 6178 9596 6184 9648
rect 6236 9596 6242 9648
rect 10042 9596 10048 9648
rect 10100 9636 10106 9648
rect 10100 9608 17264 9636
rect 10100 9596 10106 9608
rect 17126 9568 17132 9580
rect 7300 9540 17132 9568
rect 7300 9240 7328 9540
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17236 9568 17264 9608
rect 17770 9596 17776 9648
rect 17828 9636 17834 9648
rect 19978 9636 19984 9648
rect 17828 9608 19984 9636
rect 17828 9596 17834 9608
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 22186 9596 22192 9648
rect 22244 9636 22250 9648
rect 24118 9636 24124 9648
rect 22244 9608 24124 9636
rect 22244 9596 22250 9608
rect 24118 9596 24124 9608
rect 24176 9596 24182 9648
rect 28966 9636 28994 9676
rect 29270 9664 29276 9676
rect 29328 9664 29334 9716
rect 24596 9608 28994 9636
rect 29380 9636 29408 9812
rect 31726 9704 31754 9880
rect 34330 9704 34336 9716
rect 31726 9676 34336 9704
rect 34330 9664 34336 9676
rect 34388 9664 34394 9716
rect 37642 9636 37648 9648
rect 29380 9608 37648 9636
rect 23474 9568 23480 9580
rect 17236 9540 23480 9568
rect 23474 9528 23480 9540
rect 23532 9528 23538 9580
rect 23566 9528 23572 9580
rect 23624 9568 23630 9580
rect 24394 9568 24400 9580
rect 23624 9540 24400 9568
rect 23624 9528 23630 9540
rect 24394 9528 24400 9540
rect 24452 9528 24458 9580
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 21818 9500 21824 9512
rect 18656 9472 21824 9500
rect 18656 9460 18662 9472
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 24596 9500 24624 9608
rect 37642 9596 37648 9608
rect 37700 9596 37706 9648
rect 24670 9528 24676 9580
rect 24728 9568 24734 9580
rect 24728 9540 27016 9568
rect 24728 9528 24734 9540
rect 22060 9472 24624 9500
rect 22060 9460 22066 9472
rect 24762 9460 24768 9512
rect 24820 9500 24826 9512
rect 26988 9500 27016 9540
rect 28166 9528 28172 9580
rect 28224 9568 28230 9580
rect 33226 9568 33232 9580
rect 28224 9540 33232 9568
rect 28224 9528 28230 9540
rect 33226 9528 33232 9540
rect 33284 9528 33290 9580
rect 33594 9500 33600 9512
rect 24820 9472 26924 9500
rect 26988 9472 33600 9500
rect 24820 9460 24826 9472
rect 12710 9432 12716 9444
rect 7392 9404 12716 9432
rect 7282 9188 7288 9240
rect 7340 9188 7346 9240
rect 1964 9132 2774 9160
rect 1964 8832 1992 9132
rect 2746 9024 2774 9132
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 7392 9160 7420 9404
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 17402 9432 17408 9444
rect 12860 9404 17408 9432
rect 12860 9392 12866 9404
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 26510 9432 26516 9444
rect 22572 9404 26516 9432
rect 22572 9364 22600 9404
rect 26510 9392 26516 9404
rect 26568 9392 26574 9444
rect 26896 9432 26924 9472
rect 33594 9460 33600 9472
rect 33652 9460 33658 9512
rect 26896 9404 28994 9432
rect 13556 9336 22600 9364
rect 13556 9296 13584 9336
rect 24854 9324 24860 9376
rect 24912 9364 24918 9376
rect 27798 9364 27804 9376
rect 24912 9336 27804 9364
rect 24912 9324 24918 9336
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 28966 9364 28994 9404
rect 32582 9364 32588 9376
rect 28966 9336 32588 9364
rect 32582 9324 32588 9336
rect 32640 9324 32646 9376
rect 33870 9324 33876 9376
rect 33928 9364 33934 9376
rect 43806 9364 43812 9376
rect 33928 9336 43812 9364
rect 33928 9324 33934 9336
rect 43806 9324 43812 9336
rect 43864 9324 43870 9376
rect 5408 9132 7420 9160
rect 7484 9268 13584 9296
rect 5408 9120 5414 9132
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 7484 9092 7512 9268
rect 13630 9256 13636 9308
rect 13688 9296 13694 9308
rect 22370 9296 22376 9308
rect 13688 9268 22376 9296
rect 13688 9256 13694 9268
rect 22370 9256 22376 9268
rect 22428 9256 22434 9308
rect 28350 9256 28356 9308
rect 28408 9296 28414 9308
rect 34054 9296 34060 9308
rect 28408 9268 34060 9296
rect 28408 9256 28414 9268
rect 34054 9256 34060 9268
rect 34112 9256 34118 9308
rect 34606 9256 34612 9308
rect 34664 9296 34670 9308
rect 42794 9296 42800 9308
rect 34664 9268 42800 9296
rect 34664 9256 34670 9268
rect 42794 9256 42800 9268
rect 42852 9256 42858 9308
rect 9122 9188 9128 9240
rect 9180 9228 9186 9240
rect 21358 9228 21364 9240
rect 9180 9200 21364 9228
rect 9180 9188 9186 9200
rect 21358 9188 21364 9200
rect 21416 9188 21422 9240
rect 21450 9188 21456 9240
rect 21508 9228 21514 9240
rect 22186 9228 22192 9240
rect 21508 9200 22192 9228
rect 21508 9188 21514 9200
rect 22186 9188 22192 9200
rect 22244 9188 22250 9240
rect 26878 9228 26884 9240
rect 22296 9200 26884 9228
rect 11974 9160 11980 9172
rect 5040 9064 7512 9092
rect 7576 9132 11980 9160
rect 5040 9052 5046 9064
rect 7576 9024 7604 9132
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12066 9120 12072 9172
rect 12124 9160 12130 9172
rect 21634 9160 21640 9172
rect 12124 9132 21640 9160
rect 12124 9120 12130 9132
rect 21634 9120 21640 9132
rect 21692 9120 21698 9172
rect 12268 9064 14780 9092
rect 2746 8996 7604 9024
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 12268 9024 12296 9064
rect 13630 9024 13636 9036
rect 10284 8996 12296 9024
rect 12406 8996 13636 9024
rect 10284 8984 10290 8996
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 12066 8956 12072 8968
rect 10560 8928 12072 8956
rect 10560 8916 10566 8928
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 12406 8888 12434 8996
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 14752 9024 14780 9064
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 20346 9092 20352 9104
rect 17276 9064 20352 9092
rect 17276 9052 17282 9064
rect 20346 9052 20352 9064
rect 20404 9052 20410 9104
rect 22296 9092 22324 9200
rect 26878 9188 26884 9200
rect 26936 9188 26942 9240
rect 28442 9188 28448 9240
rect 28500 9228 28506 9240
rect 39114 9228 39120 9240
rect 28500 9200 39120 9228
rect 28500 9188 28506 9200
rect 39114 9188 39120 9200
rect 39172 9188 39178 9240
rect 27982 9120 27988 9172
rect 28040 9160 28046 9172
rect 33962 9160 33968 9172
rect 28040 9132 33968 9160
rect 28040 9120 28046 9132
rect 33962 9120 33968 9132
rect 34020 9120 34026 9172
rect 34330 9120 34336 9172
rect 34388 9160 34394 9172
rect 36446 9160 36452 9172
rect 34388 9132 36452 9160
rect 34388 9120 34394 9132
rect 36446 9120 36452 9132
rect 36504 9120 36510 9172
rect 22112 9064 22324 9092
rect 21634 9024 21640 9036
rect 14752 8996 21640 9024
rect 21634 8984 21640 8996
rect 21692 8984 21698 9036
rect 22112 8956 22140 9064
rect 22462 9052 22468 9104
rect 22520 9092 22526 9104
rect 25498 9092 25504 9104
rect 22520 9064 25504 9092
rect 22520 9052 22526 9064
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 29086 9052 29092 9104
rect 29144 9092 29150 9104
rect 32122 9092 32128 9104
rect 29144 9064 32128 9092
rect 29144 9052 29150 9064
rect 32122 9052 32128 9064
rect 32180 9052 32186 9104
rect 36630 9052 36636 9104
rect 36688 9092 36694 9104
rect 45462 9092 45468 9104
rect 36688 9064 45468 9092
rect 36688 9052 36694 9064
rect 45462 9052 45468 9064
rect 45520 9052 45526 9104
rect 22738 8984 22744 9036
rect 22796 9024 22802 9036
rect 24670 9024 24676 9036
rect 22796 8996 24676 9024
rect 22796 8984 22802 8996
rect 24670 8984 24676 8996
rect 24728 8984 24734 9036
rect 36538 9024 36544 9036
rect 24872 8996 36544 9024
rect 13372 8928 22140 8956
rect 13372 8900 13400 8928
rect 23106 8916 23112 8968
rect 23164 8956 23170 8968
rect 24872 8956 24900 8996
rect 36538 8984 36544 8996
rect 36596 8984 36602 9036
rect 36814 8984 36820 9036
rect 36872 9024 36878 9036
rect 45094 9024 45100 9036
rect 36872 8996 45100 9024
rect 36872 8984 36878 8996
rect 45094 8984 45100 8996
rect 45152 8984 45158 9036
rect 23164 8928 24900 8956
rect 23164 8916 23170 8928
rect 28350 8916 28356 8968
rect 28408 8956 28414 8968
rect 36998 8956 37004 8968
rect 28408 8928 37004 8956
rect 28408 8916 28414 8928
rect 36998 8916 37004 8928
rect 37056 8916 37062 8968
rect 8536 8860 12434 8888
rect 8536 8848 8542 8860
rect 13354 8848 13360 8900
rect 13412 8848 13418 8900
rect 13538 8848 13544 8900
rect 13596 8888 13602 8900
rect 22002 8888 22008 8900
rect 13596 8860 22008 8888
rect 13596 8848 13602 8860
rect 22002 8848 22008 8860
rect 22060 8848 22066 8900
rect 22462 8848 22468 8900
rect 22520 8888 22526 8900
rect 24854 8888 24860 8900
rect 22520 8860 24860 8888
rect 22520 8848 22526 8860
rect 24854 8848 24860 8860
rect 24912 8848 24918 8900
rect 36170 8888 36176 8900
rect 28092 8860 36176 8888
rect 1946 8780 1952 8832
rect 2004 8780 2010 8832
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 9674 8820 9680 8832
rect 4764 8792 9680 8820
rect 4764 8780 4770 8792
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 23014 8820 23020 8832
rect 10652 8792 23020 8820
rect 10652 8780 10658 8792
rect 23014 8780 23020 8792
rect 23072 8780 23078 8832
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 27614 8820 27620 8832
rect 24176 8792 27620 8820
rect 24176 8780 24182 8792
rect 27614 8780 27620 8792
rect 27672 8780 27678 8832
rect 27798 8780 27804 8832
rect 27856 8820 27862 8832
rect 28092 8820 28120 8860
rect 36170 8848 36176 8860
rect 36228 8848 36234 8900
rect 36262 8848 36268 8900
rect 36320 8888 36326 8900
rect 43622 8888 43628 8900
rect 36320 8860 43628 8888
rect 36320 8848 36326 8860
rect 43622 8848 43628 8860
rect 43680 8848 43686 8900
rect 27856 8792 28120 8820
rect 27856 8780 27862 8792
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 40678 8820 40684 8832
rect 34572 8792 40684 8820
rect 34572 8780 34578 8792
rect 40678 8780 40684 8792
rect 40736 8780 40742 8832
rect 1104 8730 46984 8752
rect 1104 8678 12380 8730
rect 12432 8678 12444 8730
rect 12496 8678 12508 8730
rect 12560 8678 12572 8730
rect 12624 8678 12636 8730
rect 12688 8678 23810 8730
rect 23862 8678 23874 8730
rect 23926 8678 23938 8730
rect 23990 8678 24002 8730
rect 24054 8678 24066 8730
rect 24118 8678 35240 8730
rect 35292 8678 35304 8730
rect 35356 8678 35368 8730
rect 35420 8678 35432 8730
rect 35484 8678 35496 8730
rect 35548 8678 46670 8730
rect 46722 8678 46734 8730
rect 46786 8678 46798 8730
rect 46850 8678 46862 8730
rect 46914 8678 46926 8730
rect 46978 8678 46984 8730
rect 1104 8656 46984 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2222 8616 2228 8628
rect 1811 8588 2228 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 2685 8619 2743 8625
rect 2685 8585 2697 8619
rect 2731 8616 2743 8619
rect 2958 8616 2964 8628
rect 2731 8588 2964 8616
rect 2731 8585 2743 8588
rect 2685 8579 2743 8585
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 3053 8619 3111 8625
rect 3053 8585 3065 8619
rect 3099 8616 3111 8619
rect 3326 8616 3332 8628
rect 3099 8588 3332 8616
rect 3099 8585 3111 8588
rect 3053 8579 3111 8585
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3694 8616 3700 8628
rect 3467 8588 3700 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 3973 8619 4031 8625
rect 3973 8585 3985 8619
rect 4019 8616 4031 8619
rect 4430 8616 4436 8628
rect 4019 8588 4436 8616
rect 4019 8585 4031 8588
rect 3973 8579 4031 8585
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4890 8616 4896 8628
rect 4571 8588 4896 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 4982 8576 4988 8628
rect 5040 8576 5046 8628
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5442 8616 5448 8628
rect 5123 8588 5448 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5902 8616 5908 8628
rect 5675 8588 5908 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6270 8616 6276 8628
rect 6043 8588 6276 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6730 8576 6736 8628
rect 6788 8576 6794 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7742 8616 7748 8628
rect 7147 8588 7748 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8021 8619 8079 8625
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 8202 8616 8208 8628
rect 8067 8588 8208 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 8478 8576 8484 8628
rect 8536 8576 8542 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8585 8631 8619
rect 8573 8579 8631 8585
rect 2777 8551 2835 8557
rect 2777 8517 2789 8551
rect 2823 8548 2835 8551
rect 5000 8548 5028 8576
rect 2823 8520 5028 8548
rect 5169 8551 5227 8557
rect 2823 8517 2835 8520
rect 2777 8511 2835 8517
rect 5169 8517 5181 8551
rect 5215 8548 5227 8551
rect 5350 8548 5356 8560
rect 5215 8520 5356 8548
rect 5215 8517 5227 8520
rect 5169 8511 5227 8517
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 5721 8551 5779 8557
rect 5721 8517 5733 8551
rect 5767 8548 5779 8551
rect 8496 8548 8524 8576
rect 5767 8520 8524 8548
rect 8588 8548 8616 8579
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8904 8588 9045 8616
rect 8904 8576 8910 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9490 8616 9496 8628
rect 9033 8579 9091 8585
rect 9140 8588 9496 8616
rect 9140 8548 9168 8588
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10410 8616 10416 8628
rect 10091 8588 10416 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10597 8619 10655 8625
rect 10597 8585 10609 8619
rect 10643 8616 10655 8619
rect 10962 8616 10968 8628
rect 10643 8588 10968 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11422 8616 11428 8628
rect 11195 8588 11428 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 11701 8619 11759 8625
rect 11701 8585 11713 8619
rect 11747 8616 11759 8619
rect 12158 8616 12164 8628
rect 11747 8588 12164 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12250 8576 12256 8628
rect 12308 8576 12314 8628
rect 12805 8619 12863 8625
rect 12805 8585 12817 8619
rect 12851 8616 12863 8619
rect 13262 8616 13268 8628
rect 12851 8588 13268 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 13998 8616 14004 8628
rect 13771 8588 14004 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14645 8619 14703 8625
rect 14645 8585 14657 8619
rect 14691 8616 14703 8619
rect 14918 8616 14924 8628
rect 14691 8588 14924 8616
rect 14691 8585 14703 8588
rect 14645 8579 14703 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15013 8619 15071 8625
rect 15013 8585 15025 8619
rect 15059 8616 15071 8619
rect 15470 8616 15476 8628
rect 15059 8588 15476 8616
rect 15059 8585 15071 8588
rect 15013 8579 15071 8585
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 15749 8619 15807 8625
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 16206 8616 16212 8628
rect 15795 8588 16212 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16482 8616 16488 8628
rect 16347 8588 16488 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 17310 8616 17316 8628
rect 17083 8588 17316 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 17589 8619 17647 8625
rect 17589 8585 17601 8619
rect 17635 8616 17647 8619
rect 17678 8616 17684 8628
rect 17635 8588 17684 8616
rect 17635 8585 17647 8588
rect 17589 8579 17647 8585
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 18046 8576 18052 8628
rect 18104 8576 18110 8628
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 18601 8619 18659 8625
rect 18601 8616 18613 8619
rect 18472 8588 18613 8616
rect 18472 8576 18478 8588
rect 18601 8585 18613 8588
rect 18647 8585 18659 8619
rect 18601 8579 18659 8585
rect 18782 8576 18788 8628
rect 18840 8616 18846 8628
rect 18969 8619 19027 8625
rect 18969 8616 18981 8619
rect 18840 8588 18981 8616
rect 18840 8576 18846 8588
rect 18969 8585 18981 8588
rect 19015 8585 19027 8619
rect 18969 8579 19027 8585
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 20165 8619 20223 8625
rect 20165 8616 20177 8619
rect 19944 8588 20177 8616
rect 19944 8576 19950 8588
rect 20165 8585 20177 8588
rect 20211 8585 20223 8619
rect 20165 8579 20223 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20530 8616 20536 8628
rect 20404 8588 20536 8616
rect 20404 8576 20410 8588
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 21450 8616 21456 8628
rect 21284 8588 21456 8616
rect 8588 8520 9168 8548
rect 9401 8551 9459 8557
rect 5767 8517 5779 8520
rect 5721 8511 5779 8517
rect 9401 8517 9413 8551
rect 9447 8548 9459 8551
rect 9582 8548 9588 8560
rect 9447 8520 9588 8548
rect 9447 8517 9459 8520
rect 9401 8511 9459 8517
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 9769 8551 9827 8557
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 10502 8548 10508 8560
rect 9815 8520 10508 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 10689 8551 10747 8557
rect 10689 8517 10701 8551
rect 10735 8548 10747 8551
rect 14826 8548 14832 8560
rect 10735 8520 14832 8548
rect 10735 8517 10747 8520
rect 10689 8511 10747 8517
rect 14826 8508 14832 8520
rect 14884 8508 14890 8560
rect 17126 8548 17132 8560
rect 15212 8520 17132 8548
rect 1946 8440 1952 8492
rect 2004 8440 2010 8492
rect 2314 8440 2320 8492
rect 2372 8440 2378 8492
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 2590 8412 2596 8424
rect 2148 8384 2596 8412
rect 2148 8353 2176 8384
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8313 2191 8347
rect 3620 8344 3648 8443
rect 4264 8412 4292 8443
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7190 8480 7196 8492
rect 6871 8452 7196 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 8113 8483 8171 8489
rect 7699 8452 8064 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 7926 8412 7932 8424
rect 4264 8384 7932 8412
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 6454 8344 6460 8356
rect 3620 8316 6460 8344
rect 2133 8307 2191 8313
rect 6454 8304 6460 8316
rect 6512 8304 6518 8356
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 7834 8344 7840 8356
rect 7515 8316 7840 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 7834 8304 7840 8316
rect 7892 8304 7898 8356
rect 8036 8276 8064 8452
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 9122 8480 9128 8492
rect 8711 8452 9128 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 8128 8412 8156 8443
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 10042 8480 10048 8492
rect 9263 8452 10048 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10594 8440 10600 8492
rect 10652 8440 10658 8492
rect 11241 8483 11299 8489
rect 11241 8449 11253 8483
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 10612 8412 10640 8440
rect 8128 8384 10640 8412
rect 11256 8412 11284 8443
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12802 8480 12808 8492
rect 12391 8452 12808 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8480 13875 8483
rect 14642 8480 14648 8492
rect 13863 8452 14648 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 15212 8480 15240 8520
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 19242 8508 19248 8560
rect 19300 8508 19306 8560
rect 21284 8548 21312 8588
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 22278 8616 22284 8628
rect 22020 8588 22284 8616
rect 21726 8548 21732 8560
rect 19536 8520 21312 8548
rect 21376 8520 21732 8548
rect 14783 8452 15240 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 15286 8440 15292 8492
rect 15344 8440 15350 8492
rect 15945 8483 16003 8489
rect 15945 8449 15957 8483
rect 15991 8449 16003 8483
rect 15945 8443 16003 8449
rect 16393 8483 16451 8489
rect 16393 8449 16405 8483
rect 16439 8480 16451 8483
rect 17034 8480 17040 8492
rect 16439 8452 17040 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 13556 8412 13584 8440
rect 11256 8384 13584 8412
rect 15948 8412 15976 8443
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 17954 8440 17960 8492
rect 18012 8440 18018 8492
rect 18414 8440 18420 8492
rect 18472 8440 18478 8492
rect 18782 8440 18788 8492
rect 18840 8440 18846 8492
rect 19536 8480 19564 8520
rect 19260 8452 19564 8480
rect 19260 8412 19288 8452
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 19978 8440 19984 8492
rect 20036 8440 20042 8492
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 20349 8483 20407 8489
rect 20349 8480 20361 8483
rect 20220 8452 20361 8480
rect 20220 8440 20226 8452
rect 20349 8449 20361 8452
rect 20395 8449 20407 8483
rect 20349 8443 20407 8449
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 21376 8489 21404 8520
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 21637 8483 21695 8489
rect 21637 8449 21649 8483
rect 21683 8480 21695 8483
rect 21818 8480 21824 8492
rect 21683 8452 21824 8480
rect 21683 8449 21695 8452
rect 21637 8443 21695 8449
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 22020 8489 22048 8588
rect 22278 8576 22284 8588
rect 22336 8576 22342 8628
rect 22554 8576 22560 8628
rect 22612 8576 22618 8628
rect 22646 8576 22652 8628
rect 22704 8616 22710 8628
rect 22925 8619 22983 8625
rect 22925 8616 22937 8619
rect 22704 8588 22937 8616
rect 22704 8576 22710 8588
rect 22925 8585 22937 8588
rect 22971 8585 22983 8619
rect 22925 8579 22983 8585
rect 23014 8576 23020 8628
rect 23072 8616 23078 8628
rect 24029 8619 24087 8625
rect 24029 8616 24041 8619
rect 23072 8588 24041 8616
rect 23072 8576 23078 8588
rect 24029 8585 24041 8588
rect 24075 8585 24087 8619
rect 24029 8579 24087 8585
rect 25774 8576 25780 8628
rect 25832 8616 25838 8628
rect 30653 8619 30711 8625
rect 30653 8616 30665 8619
rect 25832 8588 30665 8616
rect 25832 8576 25838 8588
rect 30653 8585 30665 8588
rect 30699 8585 30711 8619
rect 30653 8579 30711 8585
rect 30742 8576 30748 8628
rect 30800 8576 30806 8628
rect 31110 8576 31116 8628
rect 31168 8616 31174 8628
rect 31757 8619 31815 8625
rect 31757 8616 31769 8619
rect 31168 8588 31769 8616
rect 31168 8576 31174 8588
rect 31757 8585 31769 8588
rect 31803 8585 31815 8619
rect 31757 8579 31815 8585
rect 32122 8576 32128 8628
rect 32180 8576 32186 8628
rect 32493 8619 32551 8625
rect 32493 8585 32505 8619
rect 32539 8585 32551 8619
rect 32493 8579 32551 8585
rect 22572 8548 22600 8576
rect 23198 8548 23204 8560
rect 22296 8520 22600 8548
rect 22848 8520 23204 8548
rect 22296 8489 22324 8520
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8480 22431 8483
rect 22554 8480 22560 8492
rect 22419 8452 22560 8480
rect 22419 8449 22431 8452
rect 22373 8443 22431 8449
rect 22554 8440 22560 8452
rect 22612 8440 22618 8492
rect 22848 8489 22876 8520
rect 23198 8508 23204 8520
rect 23256 8508 23262 8560
rect 23750 8548 23756 8560
rect 23400 8520 23756 8548
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 23106 8440 23112 8492
rect 23164 8440 23170 8492
rect 23400 8489 23428 8520
rect 23750 8508 23756 8520
rect 23808 8508 23814 8560
rect 24302 8548 24308 8560
rect 23952 8520 24308 8548
rect 23385 8483 23443 8489
rect 23385 8449 23397 8483
rect 23431 8449 23443 8483
rect 23385 8443 23443 8449
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 23842 8480 23848 8492
rect 23707 8452 23848 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 23842 8440 23848 8452
rect 23900 8440 23906 8492
rect 23952 8489 23980 8520
rect 24302 8508 24308 8520
rect 24360 8508 24366 8560
rect 27338 8508 27344 8560
rect 27396 8548 27402 8560
rect 30374 8548 30380 8560
rect 27396 8520 30380 8548
rect 27396 8508 27402 8520
rect 30374 8508 30380 8520
rect 30432 8508 30438 8560
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 24213 8483 24271 8489
rect 24213 8449 24225 8483
rect 24259 8480 24271 8483
rect 24394 8480 24400 8492
rect 24259 8452 24400 8480
rect 24259 8449 24271 8452
rect 24213 8443 24271 8449
rect 24394 8440 24400 8452
rect 24452 8440 24458 8492
rect 24581 8483 24639 8489
rect 24581 8449 24593 8483
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 15948 8384 19288 8412
rect 19518 8372 19524 8424
rect 19576 8412 19582 8424
rect 19576 8384 20576 8412
rect 19576 8372 19582 8384
rect 13173 8347 13231 8353
rect 8220 8316 9674 8344
rect 8220 8276 8248 8316
rect 8036 8248 8248 8276
rect 9646 8276 9674 8316
rect 13173 8313 13185 8347
rect 13219 8344 13231 8347
rect 13446 8344 13452 8356
rect 13219 8316 13452 8344
rect 13219 8313 13231 8316
rect 13173 8307 13231 8313
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 14458 8304 14464 8356
rect 14516 8304 14522 8356
rect 17218 8304 17224 8356
rect 17276 8344 17282 8356
rect 19702 8344 19708 8356
rect 17276 8316 19708 8344
rect 17276 8304 17282 8316
rect 19702 8304 19708 8316
rect 19760 8304 19766 8356
rect 20548 8353 20576 8384
rect 23750 8372 23756 8424
rect 23808 8372 23814 8424
rect 24596 8412 24624 8443
rect 24946 8440 24952 8492
rect 25004 8440 25010 8492
rect 25314 8440 25320 8492
rect 25372 8440 25378 8492
rect 25682 8440 25688 8492
rect 25740 8440 25746 8492
rect 26050 8440 26056 8492
rect 26108 8440 26114 8492
rect 26418 8440 26424 8492
rect 26476 8440 26482 8492
rect 26786 8440 26792 8492
rect 26844 8440 26850 8492
rect 27154 8440 27160 8492
rect 27212 8440 27218 8492
rect 27522 8440 27528 8492
rect 27580 8440 27586 8492
rect 27890 8440 27896 8492
rect 27948 8440 27954 8492
rect 28258 8440 28264 8492
rect 28316 8440 28322 8492
rect 28626 8440 28632 8492
rect 28684 8440 28690 8492
rect 28718 8440 28724 8492
rect 28776 8480 28782 8492
rect 28997 8483 29055 8489
rect 28997 8480 29009 8483
rect 28776 8452 29009 8480
rect 28776 8440 28782 8452
rect 28997 8449 29009 8452
rect 29043 8449 29055 8483
rect 28997 8443 29055 8449
rect 29362 8440 29368 8492
rect 29420 8440 29426 8492
rect 29730 8440 29736 8492
rect 29788 8440 29794 8492
rect 30098 8440 30104 8492
rect 30156 8440 30162 8492
rect 30190 8440 30196 8492
rect 30248 8480 30254 8492
rect 30469 8483 30527 8489
rect 30469 8480 30481 8483
rect 30248 8452 30481 8480
rect 30248 8440 30254 8452
rect 30469 8449 30481 8452
rect 30515 8449 30527 8483
rect 30760 8484 30788 8576
rect 30837 8484 30895 8489
rect 30760 8483 30895 8484
rect 30760 8456 30849 8483
rect 30469 8443 30527 8449
rect 30837 8449 30849 8456
rect 30883 8449 30895 8483
rect 30837 8443 30895 8449
rect 31202 8440 31208 8492
rect 31260 8440 31266 8492
rect 31570 8440 31576 8492
rect 31628 8440 31634 8492
rect 31662 8440 31668 8492
rect 31720 8480 31726 8492
rect 31941 8483 31999 8489
rect 31941 8480 31953 8483
rect 31720 8452 31953 8480
rect 31720 8440 31726 8452
rect 31941 8449 31953 8452
rect 31987 8449 31999 8483
rect 31941 8443 31999 8449
rect 32306 8440 32312 8492
rect 32364 8440 32370 8492
rect 32508 8412 32536 8579
rect 32582 8576 32588 8628
rect 32640 8576 32646 8628
rect 33226 8576 33232 8628
rect 33284 8576 33290 8628
rect 33594 8576 33600 8628
rect 33652 8576 33658 8628
rect 33962 8576 33968 8628
rect 34020 8576 34026 8628
rect 34054 8576 34060 8628
rect 34112 8616 34118 8628
rect 34701 8619 34759 8625
rect 34701 8616 34713 8619
rect 34112 8588 34713 8616
rect 34112 8576 34118 8588
rect 34701 8585 34713 8588
rect 34747 8585 34759 8619
rect 34701 8579 34759 8585
rect 35066 8576 35072 8628
rect 35124 8616 35130 8628
rect 35437 8619 35495 8625
rect 35437 8616 35449 8619
rect 35124 8588 35449 8616
rect 35124 8576 35130 8588
rect 35437 8585 35449 8588
rect 35483 8585 35495 8619
rect 35437 8579 35495 8585
rect 36170 8576 36176 8628
rect 36228 8576 36234 8628
rect 36538 8576 36544 8628
rect 36596 8576 36602 8628
rect 36906 8576 36912 8628
rect 36964 8616 36970 8628
rect 38013 8619 38071 8625
rect 38013 8616 38025 8619
rect 36964 8588 38025 8616
rect 36964 8576 36970 8588
rect 38013 8585 38025 8588
rect 38059 8585 38071 8619
rect 38013 8579 38071 8585
rect 39114 8576 39120 8628
rect 39172 8576 39178 8628
rect 39390 8576 39396 8628
rect 39448 8616 39454 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 39448 8588 40049 8616
rect 39448 8576 39454 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 40589 8619 40647 8625
rect 40589 8585 40601 8619
rect 40635 8585 40647 8619
rect 40589 8579 40647 8585
rect 24596 8384 32536 8412
rect 32600 8412 32628 8576
rect 39758 8508 39764 8560
rect 39816 8548 39822 8560
rect 40604 8548 40632 8579
rect 40678 8576 40684 8628
rect 40736 8576 40742 8628
rect 40862 8576 40868 8628
rect 40920 8616 40926 8628
rect 41509 8619 41567 8625
rect 41509 8616 41521 8619
rect 40920 8588 41521 8616
rect 40920 8576 40926 8588
rect 41509 8585 41521 8588
rect 41555 8585 41567 8619
rect 41509 8579 41567 8585
rect 42613 8619 42671 8625
rect 42613 8585 42625 8619
rect 42659 8585 42671 8619
rect 42613 8579 42671 8585
rect 39816 8520 40632 8548
rect 40696 8548 40724 8576
rect 40696 8520 41092 8548
rect 39816 8508 39822 8520
rect 32674 8440 32680 8492
rect 32732 8440 32738 8492
rect 33042 8440 33048 8492
rect 33100 8440 33106 8492
rect 33410 8440 33416 8492
rect 33468 8440 33474 8492
rect 33778 8440 33784 8492
rect 33836 8440 33842 8492
rect 34146 8440 34152 8492
rect 34204 8440 34210 8492
rect 34238 8440 34244 8492
rect 34296 8480 34302 8492
rect 34517 8483 34575 8489
rect 34517 8480 34529 8483
rect 34296 8452 34529 8480
rect 34296 8440 34302 8452
rect 34517 8449 34529 8452
rect 34563 8449 34575 8483
rect 34517 8443 34575 8449
rect 34882 8440 34888 8492
rect 34940 8440 34946 8492
rect 34974 8440 34980 8492
rect 35032 8480 35038 8492
rect 35253 8483 35311 8489
rect 35253 8480 35265 8483
rect 35032 8452 35265 8480
rect 35032 8440 35038 8452
rect 35253 8449 35265 8452
rect 35299 8449 35311 8483
rect 35253 8443 35311 8449
rect 35618 8440 35624 8492
rect 35676 8440 35682 8492
rect 35710 8440 35716 8492
rect 35768 8480 35774 8492
rect 35989 8483 36047 8489
rect 35989 8480 36001 8483
rect 35768 8452 36001 8480
rect 35768 8440 35774 8452
rect 35989 8449 36001 8452
rect 36035 8449 36047 8483
rect 35989 8443 36047 8449
rect 36354 8440 36360 8492
rect 36412 8440 36418 8492
rect 36722 8440 36728 8492
rect 36780 8440 36786 8492
rect 37090 8440 37096 8492
rect 37148 8440 37154 8492
rect 37182 8440 37188 8492
rect 37240 8480 37246 8492
rect 37461 8483 37519 8489
rect 37461 8480 37473 8483
rect 37240 8452 37473 8480
rect 37240 8440 37246 8452
rect 37461 8449 37473 8452
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 37826 8440 37832 8492
rect 37884 8440 37890 8492
rect 38194 8440 38200 8492
rect 38252 8440 38258 8492
rect 38562 8440 38568 8492
rect 38620 8440 38626 8492
rect 38930 8440 38936 8492
rect 38988 8440 38994 8492
rect 39298 8440 39304 8492
rect 39356 8440 39362 8492
rect 39942 8440 39948 8492
rect 40000 8440 40006 8492
rect 40218 8440 40224 8492
rect 40276 8480 40282 8492
rect 40497 8483 40555 8489
rect 40497 8480 40509 8483
rect 40276 8452 40509 8480
rect 40276 8440 40282 8452
rect 40497 8449 40509 8452
rect 40543 8449 40555 8483
rect 40497 8443 40555 8449
rect 40586 8440 40592 8492
rect 40644 8480 40650 8492
rect 40957 8483 41015 8489
rect 40957 8480 40969 8483
rect 40644 8452 40969 8480
rect 40644 8440 40650 8452
rect 40957 8449 40969 8452
rect 41003 8449 41015 8483
rect 41064 8480 41092 8520
rect 41230 8508 41236 8560
rect 41288 8548 41294 8560
rect 42628 8548 42656 8579
rect 42702 8576 42708 8628
rect 42760 8616 42766 8628
rect 44269 8619 44327 8625
rect 44269 8616 44281 8619
rect 42760 8588 44281 8616
rect 42760 8576 42766 8588
rect 44269 8585 44281 8588
rect 44315 8585 44327 8619
rect 44269 8579 44327 8585
rect 44450 8576 44456 8628
rect 44508 8616 44514 8628
rect 45741 8619 45799 8625
rect 45741 8616 45753 8619
rect 44508 8588 45753 8616
rect 44508 8576 44514 8588
rect 45741 8585 45753 8588
rect 45787 8585 45799 8619
rect 45741 8579 45799 8585
rect 41288 8520 42656 8548
rect 41288 8508 41294 8520
rect 42794 8508 42800 8560
rect 42852 8548 42858 8560
rect 43073 8551 43131 8557
rect 43073 8548 43085 8551
rect 42852 8520 43085 8548
rect 42852 8508 42858 8520
rect 43073 8517 43085 8520
rect 43119 8517 43131 8551
rect 43073 8511 43131 8517
rect 43346 8508 43352 8560
rect 43404 8548 43410 8560
rect 43404 8520 45416 8548
rect 43404 8508 43410 8520
rect 41417 8483 41475 8489
rect 41417 8480 41429 8483
rect 41064 8452 41429 8480
rect 40957 8443 41015 8449
rect 41417 8449 41429 8452
rect 41463 8449 41475 8483
rect 42521 8483 42579 8489
rect 42521 8480 42533 8483
rect 41417 8443 41475 8449
rect 41524 8452 42533 8480
rect 32600 8384 32996 8412
rect 20533 8347 20591 8353
rect 20533 8313 20545 8347
rect 20579 8313 20591 8347
rect 20533 8307 20591 8313
rect 22278 8304 22284 8356
rect 22336 8344 22342 8356
rect 23477 8347 23535 8353
rect 23477 8344 23489 8347
rect 22336 8316 23489 8344
rect 22336 8304 22342 8316
rect 23477 8313 23489 8316
rect 23523 8313 23535 8347
rect 23768 8344 23796 8372
rect 24397 8347 24455 8353
rect 24397 8344 24409 8347
rect 23768 8316 24409 8344
rect 23477 8307 23535 8313
rect 24397 8313 24409 8316
rect 24443 8313 24455 8347
rect 24397 8307 24455 8313
rect 26142 8304 26148 8356
rect 26200 8344 26206 8356
rect 26237 8347 26295 8353
rect 26237 8344 26249 8347
rect 26200 8316 26249 8344
rect 26200 8304 26206 8316
rect 26237 8313 26249 8316
rect 26283 8313 26295 8347
rect 26237 8307 26295 8313
rect 27430 8304 27436 8356
rect 27488 8344 27494 8356
rect 27709 8347 27767 8353
rect 27709 8344 27721 8347
rect 27488 8316 27721 8344
rect 27488 8304 27494 8316
rect 27709 8313 27721 8316
rect 27755 8313 27767 8347
rect 28077 8347 28135 8353
rect 28077 8344 28089 8347
rect 27709 8307 27767 8313
rect 27816 8316 28089 8344
rect 14476 8276 14504 8304
rect 9646 8248 14504 8276
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 20901 8279 20959 8285
rect 20901 8276 20913 8279
rect 20772 8248 20913 8276
rect 20772 8236 20778 8248
rect 20901 8245 20913 8248
rect 20947 8245 20959 8279
rect 20901 8239 20959 8245
rect 21174 8236 21180 8288
rect 21232 8236 21238 8288
rect 21450 8236 21456 8288
rect 21508 8236 21514 8288
rect 21818 8236 21824 8288
rect 21876 8236 21882 8288
rect 22002 8236 22008 8288
rect 22060 8276 22066 8288
rect 22097 8279 22155 8285
rect 22097 8276 22109 8279
rect 22060 8248 22109 8276
rect 22060 8236 22066 8248
rect 22097 8245 22109 8248
rect 22143 8245 22155 8279
rect 22097 8239 22155 8245
rect 22554 8236 22560 8288
rect 22612 8236 22618 8288
rect 22646 8236 22652 8288
rect 22704 8236 22710 8288
rect 22738 8236 22744 8288
rect 22796 8276 22802 8288
rect 23201 8279 23259 8285
rect 23201 8276 23213 8279
rect 22796 8248 23213 8276
rect 22796 8236 22802 8248
rect 23201 8245 23213 8248
rect 23247 8245 23259 8279
rect 23201 8239 23259 8245
rect 23566 8236 23572 8288
rect 23624 8276 23630 8288
rect 23753 8279 23811 8285
rect 23753 8276 23765 8279
rect 23624 8248 23765 8276
rect 23624 8236 23630 8248
rect 23753 8245 23765 8248
rect 23799 8245 23811 8279
rect 23753 8239 23811 8245
rect 24762 8236 24768 8288
rect 24820 8236 24826 8288
rect 25130 8236 25136 8288
rect 25188 8236 25194 8288
rect 25222 8236 25228 8288
rect 25280 8276 25286 8288
rect 25501 8279 25559 8285
rect 25501 8276 25513 8279
rect 25280 8248 25513 8276
rect 25280 8236 25286 8248
rect 25501 8245 25513 8248
rect 25547 8245 25559 8279
rect 25501 8239 25559 8245
rect 25866 8236 25872 8288
rect 25924 8236 25930 8288
rect 26602 8236 26608 8288
rect 26660 8236 26666 8288
rect 26786 8236 26792 8288
rect 26844 8276 26850 8288
rect 26973 8279 27031 8285
rect 26973 8276 26985 8279
rect 26844 8248 26985 8276
rect 26844 8236 26850 8248
rect 26973 8245 26985 8248
rect 27019 8245 27031 8279
rect 26973 8239 27031 8245
rect 27154 8236 27160 8288
rect 27212 8276 27218 8288
rect 27341 8279 27399 8285
rect 27341 8276 27353 8279
rect 27212 8248 27353 8276
rect 27212 8236 27218 8248
rect 27341 8245 27353 8248
rect 27387 8245 27399 8279
rect 27341 8239 27399 8245
rect 27522 8236 27528 8288
rect 27580 8276 27586 8288
rect 27816 8276 27844 8316
rect 28077 8313 28089 8316
rect 28123 8313 28135 8347
rect 28077 8307 28135 8313
rect 28994 8304 29000 8356
rect 29052 8344 29058 8356
rect 32861 8347 32919 8353
rect 32861 8344 32873 8347
rect 29052 8316 32873 8344
rect 29052 8304 29058 8316
rect 32861 8313 32873 8316
rect 32907 8313 32919 8347
rect 32968 8344 32996 8384
rect 33686 8372 33692 8424
rect 33744 8412 33750 8424
rect 41524 8412 41552 8452
rect 42521 8449 42533 8452
rect 42567 8449 42579 8483
rect 42521 8443 42579 8449
rect 43622 8440 43628 8492
rect 43680 8440 43686 8492
rect 43806 8440 43812 8492
rect 43864 8480 43870 8492
rect 44177 8483 44235 8489
rect 44177 8480 44189 8483
rect 43864 8452 44189 8480
rect 43864 8440 43870 8452
rect 44177 8449 44189 8452
rect 44223 8449 44235 8483
rect 44177 8443 44235 8449
rect 45094 8440 45100 8492
rect 45152 8440 45158 8492
rect 33744 8384 41552 8412
rect 33744 8372 33750 8384
rect 41966 8372 41972 8424
rect 42024 8412 42030 8424
rect 45388 8421 45416 8520
rect 45462 8508 45468 8560
rect 45520 8548 45526 8560
rect 45649 8551 45707 8557
rect 45649 8548 45661 8551
rect 45520 8520 45661 8548
rect 45520 8508 45526 8520
rect 45649 8517 45661 8520
rect 45695 8517 45707 8551
rect 45649 8511 45707 8517
rect 45373 8415 45431 8421
rect 42024 8384 43852 8412
rect 42024 8372 42030 8384
rect 34333 8347 34391 8353
rect 34333 8344 34345 8347
rect 32968 8316 34345 8344
rect 32861 8307 32919 8313
rect 34333 8313 34345 8316
rect 34379 8313 34391 8347
rect 34333 8307 34391 8313
rect 35066 8304 35072 8356
rect 35124 8304 35130 8356
rect 35802 8304 35808 8356
rect 35860 8304 35866 8356
rect 36446 8304 36452 8356
rect 36504 8344 36510 8356
rect 36909 8347 36967 8353
rect 36909 8344 36921 8347
rect 36504 8316 36921 8344
rect 36504 8304 36510 8316
rect 36909 8313 36921 8316
rect 36955 8313 36967 8347
rect 36909 8307 36967 8313
rect 36998 8304 37004 8356
rect 37056 8304 37062 8356
rect 37090 8304 37096 8356
rect 37148 8344 37154 8356
rect 38381 8347 38439 8353
rect 38381 8344 38393 8347
rect 37148 8316 38393 8344
rect 37148 8304 37154 8316
rect 38381 8313 38393 8316
rect 38427 8313 38439 8347
rect 38381 8307 38439 8313
rect 38746 8304 38752 8356
rect 38804 8304 38810 8356
rect 40126 8304 40132 8356
rect 40184 8344 40190 8356
rect 41141 8347 41199 8353
rect 41141 8344 41153 8347
rect 40184 8316 41153 8344
rect 40184 8304 40190 8316
rect 41141 8313 41153 8316
rect 41187 8313 41199 8347
rect 41141 8307 41199 8313
rect 41598 8304 41604 8356
rect 41656 8344 41662 8356
rect 43824 8353 43852 8384
rect 45373 8381 45385 8415
rect 45419 8381 45431 8415
rect 45373 8375 45431 8381
rect 43257 8347 43315 8353
rect 43257 8344 43269 8347
rect 41656 8316 43269 8344
rect 41656 8304 41662 8316
rect 43257 8313 43269 8316
rect 43303 8313 43315 8347
rect 43257 8307 43315 8313
rect 43809 8347 43867 8353
rect 43809 8313 43821 8347
rect 43855 8313 43867 8347
rect 43809 8307 43867 8313
rect 27580 8248 27844 8276
rect 27580 8236 27586 8248
rect 28166 8236 28172 8288
rect 28224 8276 28230 8288
rect 28445 8279 28503 8285
rect 28445 8276 28457 8279
rect 28224 8248 28457 8276
rect 28224 8236 28230 8248
rect 28445 8245 28457 8248
rect 28491 8245 28503 8279
rect 28445 8239 28503 8245
rect 28534 8236 28540 8288
rect 28592 8276 28598 8288
rect 28813 8279 28871 8285
rect 28813 8276 28825 8279
rect 28592 8248 28825 8276
rect 28592 8236 28598 8248
rect 28813 8245 28825 8248
rect 28859 8245 28871 8279
rect 28813 8239 28871 8245
rect 29178 8236 29184 8288
rect 29236 8236 29242 8288
rect 29270 8236 29276 8288
rect 29328 8276 29334 8288
rect 29549 8279 29607 8285
rect 29549 8276 29561 8279
rect 29328 8248 29561 8276
rect 29328 8236 29334 8248
rect 29549 8245 29561 8248
rect 29595 8245 29607 8279
rect 29549 8239 29607 8245
rect 29914 8236 29920 8288
rect 29972 8236 29978 8288
rect 30282 8236 30288 8288
rect 30340 8236 30346 8288
rect 30374 8236 30380 8288
rect 30432 8276 30438 8288
rect 31021 8279 31079 8285
rect 31021 8276 31033 8279
rect 30432 8248 31033 8276
rect 30432 8236 30438 8248
rect 31021 8245 31033 8248
rect 31067 8245 31079 8279
rect 31021 8239 31079 8245
rect 31386 8236 31392 8288
rect 31444 8236 31450 8288
rect 37016 8276 37044 8304
rect 37277 8279 37335 8285
rect 37277 8276 37289 8279
rect 37016 8248 37289 8276
rect 37277 8245 37289 8248
rect 37323 8245 37335 8279
rect 37277 8239 37335 8245
rect 37642 8236 37648 8288
rect 37700 8236 37706 8288
rect 1104 8186 46828 8208
rect 1104 8134 6665 8186
rect 6717 8134 6729 8186
rect 6781 8134 6793 8186
rect 6845 8134 6857 8186
rect 6909 8134 6921 8186
rect 6973 8134 18095 8186
rect 18147 8134 18159 8186
rect 18211 8134 18223 8186
rect 18275 8134 18287 8186
rect 18339 8134 18351 8186
rect 18403 8134 29525 8186
rect 29577 8134 29589 8186
rect 29641 8134 29653 8186
rect 29705 8134 29717 8186
rect 29769 8134 29781 8186
rect 29833 8134 40955 8186
rect 41007 8134 41019 8186
rect 41071 8134 41083 8186
rect 41135 8134 41147 8186
rect 41199 8134 41211 8186
rect 41263 8134 46828 8186
rect 1104 8112 46828 8134
rect 1118 8032 1124 8084
rect 1176 8072 1182 8084
rect 1857 8075 1915 8081
rect 1857 8072 1869 8075
rect 1176 8044 1869 8072
rect 1176 8032 1182 8044
rect 1857 8041 1869 8044
rect 1903 8041 1915 8075
rect 1857 8035 1915 8041
rect 4062 8032 4068 8084
rect 4120 8032 4126 8084
rect 4617 8075 4675 8081
rect 4617 8041 4629 8075
rect 4663 8072 4675 8075
rect 4798 8072 4804 8084
rect 4663 8044 4804 8072
rect 4663 8041 4675 8044
rect 4617 8035 4675 8041
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6604 8044 6653 8072
rect 6604 8032 6610 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7374 8072 7380 8084
rect 7239 8044 7380 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 9214 8032 9220 8084
rect 9272 8032 9278 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10318 8072 10324 8084
rect 10091 8044 10324 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 11790 8032 11796 8084
rect 11848 8032 11854 8084
rect 12621 8075 12679 8081
rect 12621 8041 12633 8075
rect 12667 8072 12679 8075
rect 12894 8072 12900 8084
rect 12667 8044 12900 8072
rect 12667 8041 12679 8044
rect 12621 8035 12679 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 14366 8032 14372 8084
rect 14424 8032 14430 8084
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 14921 8075 14979 8081
rect 14921 8072 14933 8075
rect 14792 8044 14933 8072
rect 14792 8032 14798 8044
rect 14921 8041 14933 8044
rect 14967 8041 14979 8075
rect 14921 8035 14979 8041
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 15838 8072 15844 8084
rect 15611 8044 15844 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 16666 8072 16672 8084
rect 15948 8044 16672 8072
rect 2409 8007 2467 8013
rect 2409 7973 2421 8007
rect 2455 7973 2467 8007
rect 15948 8004 15976 8044
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 17000 8044 17049 8072
rect 17000 8032 17006 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17037 8035 17095 8041
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17736 8044 17785 8072
rect 17736 8032 17742 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 17773 8035 17831 8041
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18049 8075 18107 8081
rect 18049 8072 18061 8075
rect 18012 8044 18061 8072
rect 18012 8032 18018 8044
rect 18049 8041 18061 8044
rect 18095 8041 18107 8075
rect 18049 8035 18107 8041
rect 18325 8075 18383 8081
rect 18325 8041 18337 8075
rect 18371 8072 18383 8075
rect 18414 8072 18420 8084
rect 18371 8044 18420 8072
rect 18371 8041 18383 8044
rect 18325 8035 18383 8041
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 18782 8032 18788 8084
rect 18840 8032 18846 8084
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 19576 8044 19625 8072
rect 19576 8032 19582 8044
rect 19613 8041 19625 8044
rect 19659 8041 19671 8075
rect 19613 8035 19671 8041
rect 19889 8075 19947 8081
rect 19889 8041 19901 8075
rect 19935 8072 19947 8075
rect 19978 8072 19984 8084
rect 19935 8044 19984 8072
rect 19935 8041 19947 8044
rect 19889 8035 19947 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20441 8075 20499 8081
rect 20441 8041 20453 8075
rect 20487 8041 20499 8075
rect 20441 8035 20499 8041
rect 2409 7967 2467 7973
rect 10244 7976 15976 8004
rect 1854 7896 1860 7948
rect 1912 7936 1918 7948
rect 2424 7936 2452 7967
rect 1912 7908 2452 7936
rect 1912 7896 1918 7908
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2130 7760 2136 7812
rect 2188 7760 2194 7812
rect 2608 7732 2636 7831
rect 4798 7828 4804 7880
rect 4856 7828 4862 7880
rect 10244 7877 10272 7976
rect 16390 7964 16396 8016
rect 16448 8004 16454 8016
rect 20456 8004 20484 8035
rect 20530 8032 20536 8084
rect 20588 8072 20594 8084
rect 20717 8075 20775 8081
rect 20717 8072 20729 8075
rect 20588 8044 20729 8072
rect 20588 8032 20594 8044
rect 20717 8041 20729 8044
rect 20763 8041 20775 8075
rect 20717 8035 20775 8041
rect 20898 8032 20904 8084
rect 20956 8072 20962 8084
rect 20993 8075 21051 8081
rect 20993 8072 21005 8075
rect 20956 8044 21005 8072
rect 20956 8032 20962 8044
rect 20993 8041 21005 8044
rect 21039 8041 21051 8075
rect 20993 8035 21051 8041
rect 21266 8032 21272 8084
rect 21324 8032 21330 8084
rect 21358 8032 21364 8084
rect 21416 8072 21422 8084
rect 21821 8075 21879 8081
rect 21821 8072 21833 8075
rect 21416 8044 21833 8072
rect 21416 8032 21422 8044
rect 21821 8041 21833 8044
rect 21867 8041 21879 8075
rect 21821 8035 21879 8041
rect 22370 8032 22376 8084
rect 22428 8072 22434 8084
rect 22428 8044 22784 8072
rect 22428 8032 22434 8044
rect 22649 8007 22707 8013
rect 22649 8004 22661 8007
rect 16448 7976 20484 8004
rect 20548 7976 22661 8004
rect 16448 7964 16454 7976
rect 18138 7936 18144 7948
rect 10336 7908 18144 7936
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 10229 7871 10287 7877
rect 7423 7840 10180 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 4338 7760 4344 7812
rect 4396 7760 4402 7812
rect 6914 7760 6920 7812
rect 6972 7760 6978 7812
rect 9493 7803 9551 7809
rect 9493 7769 9505 7803
rect 9539 7800 9551 7803
rect 10042 7800 10048 7812
rect 9539 7772 10048 7800
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 10152 7800 10180 7840
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10336 7800 10364 7908
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 19702 7936 19708 7948
rect 19076 7908 19708 7936
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 13722 7868 13728 7880
rect 12851 7840 13728 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 15105 7871 15163 7877
rect 14568 7840 14872 7868
rect 10152 7772 10364 7800
rect 12069 7803 12127 7809
rect 12069 7769 12081 7803
rect 12115 7800 12127 7803
rect 14568 7800 14596 7840
rect 14844 7812 14872 7840
rect 15105 7837 15117 7871
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 12115 7772 14596 7800
rect 12115 7769 12127 7772
rect 12069 7763 12127 7769
rect 14642 7760 14648 7812
rect 14700 7760 14706 7812
rect 14826 7760 14832 7812
rect 14884 7760 14890 7812
rect 15120 7800 15148 7831
rect 15746 7828 15752 7880
rect 15804 7828 15810 7880
rect 17218 7828 17224 7880
rect 17276 7828 17282 7880
rect 17954 7828 17960 7880
rect 18012 7828 18018 7880
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18414 7868 18420 7880
rect 18279 7840 18420 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 18506 7828 18512 7880
rect 18564 7828 18570 7880
rect 18601 7871 18659 7877
rect 18601 7837 18613 7871
rect 18647 7868 18659 7871
rect 18966 7868 18972 7880
rect 18647 7840 18972 7868
rect 18647 7837 18659 7840
rect 18601 7831 18659 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19076 7877 19104 7908
rect 19702 7896 19708 7908
rect 19760 7896 19766 7948
rect 20438 7936 20444 7948
rect 19812 7908 20444 7936
rect 19061 7871 19119 7877
rect 19061 7837 19073 7871
rect 19107 7837 19119 7871
rect 19061 7831 19119 7837
rect 19518 7828 19524 7880
rect 19576 7828 19582 7880
rect 19812 7877 19840 7908
rect 20438 7896 20444 7908
rect 20496 7896 20502 7948
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 20070 7828 20076 7880
rect 20128 7828 20134 7880
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20548 7800 20576 7976
rect 22649 7973 22661 7976
rect 22695 7973 22707 8007
rect 22756 8004 22784 8044
rect 23474 8032 23480 8084
rect 23532 8072 23538 8084
rect 23753 8075 23811 8081
rect 23753 8072 23765 8075
rect 23532 8044 23765 8072
rect 23532 8032 23538 8044
rect 23753 8041 23765 8044
rect 23799 8041 23811 8075
rect 23753 8035 23811 8041
rect 24210 8032 24216 8084
rect 24268 8072 24274 8084
rect 24489 8075 24547 8081
rect 24489 8072 24501 8075
rect 24268 8044 24501 8072
rect 24268 8032 24274 8044
rect 24489 8041 24501 8044
rect 24535 8041 24547 8075
rect 24489 8035 24547 8041
rect 25130 8032 25136 8084
rect 25188 8032 25194 8084
rect 25406 8032 25412 8084
rect 25464 8032 25470 8084
rect 25498 8032 25504 8084
rect 25556 8072 25562 8084
rect 25685 8075 25743 8081
rect 25685 8072 25697 8075
rect 25556 8044 25697 8072
rect 25556 8032 25562 8044
rect 25685 8041 25697 8044
rect 25731 8041 25743 8075
rect 25685 8035 25743 8041
rect 25866 8032 25872 8084
rect 25924 8032 25930 8084
rect 27338 8072 27344 8084
rect 25976 8044 27344 8072
rect 24029 8007 24087 8013
rect 24029 8004 24041 8007
rect 22756 7976 24041 8004
rect 22649 7967 22707 7973
rect 24029 7973 24041 7976
rect 24075 7973 24087 8007
rect 25038 8004 25044 8016
rect 24029 7967 24087 7973
rect 24136 7976 25044 8004
rect 22462 7936 22468 7948
rect 20916 7908 22468 7936
rect 20625 7871 20683 7877
rect 20625 7837 20637 7871
rect 20671 7868 20683 7871
rect 20714 7868 20720 7880
rect 20671 7840 20720 7868
rect 20671 7837 20683 7840
rect 20625 7831 20683 7837
rect 20714 7828 20720 7840
rect 20772 7828 20778 7880
rect 20916 7877 20944 7908
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 22738 7936 22744 7948
rect 22572 7908 22744 7936
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21174 7828 21180 7880
rect 21232 7828 21238 7880
rect 21450 7828 21456 7880
rect 21508 7828 21514 7880
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7868 21787 7871
rect 21818 7868 21824 7880
rect 21775 7840 21824 7868
rect 21775 7837 21787 7840
rect 21729 7831 21787 7837
rect 21818 7828 21824 7840
rect 21876 7828 21882 7880
rect 22002 7828 22008 7880
rect 22060 7828 22066 7880
rect 22572 7877 22600 7908
rect 22738 7896 22744 7908
rect 22796 7896 22802 7948
rect 22281 7871 22339 7877
rect 22281 7837 22293 7871
rect 22327 7837 22339 7871
rect 22281 7831 22339 7837
rect 22557 7871 22615 7877
rect 22557 7837 22569 7871
rect 22603 7837 22615 7871
rect 22557 7831 22615 7837
rect 22296 7800 22324 7831
rect 22646 7828 22652 7880
rect 22704 7828 22710 7880
rect 22830 7828 22836 7880
rect 22888 7828 22894 7880
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23290 7868 23296 7880
rect 23155 7840 23296 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 23385 7871 23443 7877
rect 23385 7837 23397 7871
rect 23431 7868 23443 7871
rect 23566 7868 23572 7880
rect 23431 7840 23572 7868
rect 23431 7837 23443 7840
rect 23385 7831 23443 7837
rect 23566 7828 23572 7840
rect 23624 7828 23630 7880
rect 23661 7871 23719 7877
rect 23661 7837 23673 7871
rect 23707 7837 23719 7871
rect 23661 7831 23719 7837
rect 23937 7871 23995 7877
rect 23937 7837 23949 7871
rect 23983 7868 23995 7871
rect 24136 7868 24164 7976
rect 25038 7964 25044 7976
rect 25096 7964 25102 8016
rect 25148 7936 25176 8032
rect 25884 7936 25912 8032
rect 24228 7908 25176 7936
rect 25332 7908 25912 7936
rect 24228 7877 24256 7908
rect 23983 7840 24164 7868
rect 24213 7871 24271 7877
rect 23983 7837 23995 7840
rect 23937 7831 23995 7837
rect 24213 7837 24225 7871
rect 24259 7837 24271 7871
rect 24213 7831 24271 7837
rect 24673 7871 24731 7877
rect 24673 7837 24685 7871
rect 24719 7868 24731 7871
rect 24854 7868 24860 7880
rect 24719 7840 24860 7868
rect 24719 7837 24731 7840
rect 24673 7831 24731 7837
rect 22664 7800 22692 7828
rect 15120 7772 20576 7800
rect 20640 7772 22140 7800
rect 22296 7772 22692 7800
rect 20640 7744 20668 7772
rect 15102 7732 15108 7744
rect 2608 7704 15108 7732
rect 15102 7692 15108 7704
rect 15160 7692 15166 7744
rect 16206 7692 16212 7744
rect 16264 7732 16270 7744
rect 18877 7735 18935 7741
rect 18877 7732 18889 7735
rect 16264 7704 18889 7732
rect 16264 7692 16270 7704
rect 18877 7701 18889 7704
rect 18923 7701 18935 7735
rect 18877 7695 18935 7701
rect 19334 7692 19340 7744
rect 19392 7692 19398 7744
rect 19978 7692 19984 7744
rect 20036 7732 20042 7744
rect 20165 7735 20223 7741
rect 20165 7732 20177 7735
rect 20036 7704 20177 7732
rect 20036 7692 20042 7704
rect 20165 7701 20177 7704
rect 20211 7701 20223 7735
rect 20165 7695 20223 7701
rect 20622 7692 20628 7744
rect 20680 7692 20686 7744
rect 21542 7692 21548 7744
rect 21600 7692 21606 7744
rect 22112 7741 22140 7772
rect 22738 7760 22744 7812
rect 22796 7800 22802 7812
rect 23676 7800 23704 7831
rect 24854 7828 24860 7840
rect 24912 7828 24918 7880
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7868 25007 7871
rect 25222 7868 25228 7880
rect 24995 7840 25228 7868
rect 24995 7837 25007 7840
rect 24949 7831 25007 7837
rect 25222 7828 25228 7840
rect 25280 7828 25286 7880
rect 25332 7877 25360 7908
rect 25317 7871 25375 7877
rect 25317 7837 25329 7871
rect 25363 7837 25375 7871
rect 25317 7831 25375 7837
rect 25593 7871 25651 7877
rect 25593 7837 25605 7871
rect 25639 7868 25651 7871
rect 25774 7868 25780 7880
rect 25639 7840 25780 7868
rect 25639 7837 25651 7840
rect 25593 7831 25651 7837
rect 25774 7828 25780 7840
rect 25832 7828 25838 7880
rect 25869 7871 25927 7877
rect 25869 7837 25881 7871
rect 25915 7868 25927 7871
rect 25976 7868 26004 8044
rect 27338 8032 27344 8044
rect 27396 8032 27402 8084
rect 27706 8032 27712 8084
rect 27764 8032 27770 8084
rect 28074 8032 28080 8084
rect 28132 8032 28138 8084
rect 28445 8075 28503 8081
rect 28445 8041 28457 8075
rect 28491 8072 28503 8075
rect 28810 8072 28816 8084
rect 28491 8044 28816 8072
rect 28491 8041 28503 8044
rect 28445 8035 28503 8041
rect 28810 8032 28816 8044
rect 28868 8032 28874 8084
rect 29178 8032 29184 8084
rect 29236 8032 29242 8084
rect 29362 8032 29368 8084
rect 29420 8072 29426 8084
rect 29641 8075 29699 8081
rect 29641 8072 29653 8075
rect 29420 8044 29653 8072
rect 29420 8032 29426 8044
rect 29641 8041 29653 8044
rect 29687 8041 29699 8075
rect 29641 8035 29699 8041
rect 29914 8032 29920 8084
rect 29972 8032 29978 8084
rect 40494 8032 40500 8084
rect 40552 8072 40558 8084
rect 41141 8075 41199 8081
rect 41141 8072 41153 8075
rect 40552 8044 41153 8072
rect 40552 8032 40558 8044
rect 41141 8041 41153 8044
rect 41187 8041 41199 8075
rect 41141 8035 41199 8041
rect 42794 8032 42800 8084
rect 42852 8072 42858 8084
rect 43349 8075 43407 8081
rect 43349 8072 43361 8075
rect 42852 8044 43361 8072
rect 42852 8032 42858 8044
rect 43349 8041 43361 8044
rect 43395 8041 43407 8075
rect 43349 8035 43407 8041
rect 43714 8032 43720 8084
rect 43772 8072 43778 8084
rect 45189 8075 45247 8081
rect 45189 8072 45201 8075
rect 43772 8044 45201 8072
rect 43772 8032 43778 8044
rect 45189 8041 45201 8044
rect 45235 8041 45247 8075
rect 45189 8035 45247 8041
rect 45925 8075 45983 8081
rect 45925 8041 45937 8075
rect 45971 8072 45983 8075
rect 46566 8072 46572 8084
rect 45971 8044 46572 8072
rect 45971 8041 45983 8044
rect 45925 8035 45983 8041
rect 46566 8032 46572 8044
rect 46624 8032 46630 8084
rect 26510 7964 26516 8016
rect 26568 7964 26574 8016
rect 27062 7964 27068 8016
rect 27120 7964 27126 8016
rect 29196 7936 29224 8032
rect 29932 7936 29960 8032
rect 44174 7964 44180 8016
rect 44232 7964 44238 8016
rect 28644 7908 29224 7936
rect 29380 7908 29960 7936
rect 25915 7840 26004 7868
rect 25915 7837 25927 7840
rect 25869 7831 25927 7837
rect 26142 7828 26148 7880
rect 26200 7828 26206 7880
rect 26421 7871 26479 7877
rect 26421 7837 26433 7871
rect 26467 7868 26479 7871
rect 26602 7868 26608 7880
rect 26467 7840 26608 7868
rect 26467 7837 26479 7840
rect 26421 7831 26479 7837
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 26697 7871 26755 7877
rect 26697 7837 26709 7871
rect 26743 7868 26755 7871
rect 26786 7868 26792 7880
rect 26743 7840 26792 7868
rect 26743 7837 26755 7840
rect 26697 7831 26755 7837
rect 26786 7828 26792 7840
rect 26844 7828 26850 7880
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7868 27031 7871
rect 27154 7868 27160 7880
rect 27019 7840 27160 7868
rect 27019 7837 27031 7840
rect 26973 7831 27031 7837
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7868 27307 7871
rect 27430 7868 27436 7880
rect 27295 7840 27436 7868
rect 27295 7837 27307 7840
rect 27249 7831 27307 7837
rect 27430 7828 27436 7840
rect 27488 7828 27494 7880
rect 27522 7828 27528 7880
rect 27580 7828 27586 7880
rect 27893 7871 27951 7877
rect 27893 7837 27905 7871
rect 27939 7868 27951 7871
rect 28166 7868 28172 7880
rect 27939 7840 28172 7868
rect 27939 7837 27951 7840
rect 27893 7831 27951 7837
rect 28166 7828 28172 7840
rect 28224 7828 28230 7880
rect 28261 7871 28319 7877
rect 28261 7837 28273 7871
rect 28307 7868 28319 7871
rect 28534 7868 28540 7880
rect 28307 7840 28540 7868
rect 28307 7837 28319 7840
rect 28261 7831 28319 7837
rect 28534 7828 28540 7840
rect 28592 7828 28598 7880
rect 28644 7877 28672 7908
rect 28629 7871 28687 7877
rect 28629 7837 28641 7871
rect 28675 7837 28687 7871
rect 28629 7831 28687 7837
rect 28997 7871 29055 7877
rect 28997 7837 29009 7871
rect 29043 7868 29055 7871
rect 29270 7868 29276 7880
rect 29043 7840 29276 7868
rect 29043 7837 29055 7840
rect 28997 7831 29055 7837
rect 29270 7828 29276 7840
rect 29328 7828 29334 7880
rect 29380 7877 29408 7908
rect 29365 7871 29423 7877
rect 29365 7837 29377 7871
rect 29411 7837 29423 7871
rect 29365 7831 29423 7837
rect 29825 7871 29883 7877
rect 29825 7837 29837 7871
rect 29871 7868 29883 7871
rect 30282 7868 30288 7880
rect 29871 7840 30288 7868
rect 29871 7837 29883 7840
rect 29825 7831 29883 7837
rect 30282 7828 30288 7840
rect 30340 7828 30346 7880
rect 40034 7828 40040 7880
rect 40092 7868 40098 7880
rect 40957 7871 41015 7877
rect 40957 7868 40969 7871
rect 40092 7840 40969 7868
rect 40092 7828 40098 7840
rect 40957 7837 40969 7840
rect 41003 7837 41015 7871
rect 40957 7831 41015 7837
rect 37090 7800 37096 7812
rect 22796 7772 23520 7800
rect 23676 7772 37096 7800
rect 22796 7760 22802 7772
rect 22097 7735 22155 7741
rect 22097 7701 22109 7735
rect 22143 7701 22155 7735
rect 22097 7695 22155 7701
rect 22278 7692 22284 7744
rect 22336 7732 22342 7744
rect 22373 7735 22431 7741
rect 22373 7732 22385 7735
rect 22336 7704 22385 7732
rect 22336 7692 22342 7704
rect 22373 7701 22385 7704
rect 22419 7701 22431 7735
rect 22373 7695 22431 7701
rect 22922 7692 22928 7744
rect 22980 7692 22986 7744
rect 23198 7692 23204 7744
rect 23256 7692 23262 7744
rect 23492 7741 23520 7772
rect 37090 7760 37096 7772
rect 37148 7760 37154 7812
rect 43254 7760 43260 7812
rect 43312 7760 43318 7812
rect 43990 7760 43996 7812
rect 44048 7760 44054 7812
rect 45094 7760 45100 7812
rect 45152 7760 45158 7812
rect 45649 7803 45707 7809
rect 45649 7769 45661 7803
rect 45695 7800 45707 7803
rect 45830 7800 45836 7812
rect 45695 7772 45836 7800
rect 45695 7769 45707 7772
rect 45649 7763 45707 7769
rect 45830 7760 45836 7772
rect 45888 7760 45894 7812
rect 23477 7735 23535 7741
rect 23477 7701 23489 7735
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 24578 7692 24584 7744
rect 24636 7732 24642 7744
rect 24765 7735 24823 7741
rect 24765 7732 24777 7735
rect 24636 7704 24777 7732
rect 24636 7692 24642 7704
rect 24765 7701 24777 7704
rect 24811 7701 24823 7735
rect 24765 7695 24823 7701
rect 25130 7692 25136 7744
rect 25188 7692 25194 7744
rect 25958 7692 25964 7744
rect 26016 7692 26022 7744
rect 26234 7692 26240 7744
rect 26292 7692 26298 7744
rect 26786 7692 26792 7744
rect 26844 7692 26850 7744
rect 26878 7692 26884 7744
rect 26936 7732 26942 7744
rect 27341 7735 27399 7741
rect 27341 7732 27353 7735
rect 26936 7704 27353 7732
rect 26936 7692 26942 7704
rect 27341 7701 27353 7704
rect 27387 7701 27399 7735
rect 27341 7695 27399 7701
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 28813 7735 28871 7741
rect 28813 7732 28825 7735
rect 27672 7704 28825 7732
rect 27672 7692 27678 7704
rect 28813 7701 28825 7704
rect 28859 7701 28871 7735
rect 28813 7695 28871 7701
rect 29178 7692 29184 7744
rect 29236 7692 29242 7744
rect 1104 7642 46984 7664
rect 1104 7590 12380 7642
rect 12432 7590 12444 7642
rect 12496 7590 12508 7642
rect 12560 7590 12572 7642
rect 12624 7590 12636 7642
rect 12688 7590 23810 7642
rect 23862 7590 23874 7642
rect 23926 7590 23938 7642
rect 23990 7590 24002 7642
rect 24054 7590 24066 7642
rect 24118 7590 35240 7642
rect 35292 7590 35304 7642
rect 35356 7590 35368 7642
rect 35420 7590 35432 7642
rect 35484 7590 35496 7642
rect 35548 7590 46670 7642
rect 46722 7590 46734 7642
rect 46786 7590 46798 7642
rect 46850 7590 46862 7642
rect 46914 7590 46926 7642
rect 46978 7590 46984 7642
rect 1104 7568 46984 7590
rect 1486 7488 1492 7540
rect 1544 7488 1550 7540
rect 2130 7488 2136 7540
rect 2188 7488 2194 7540
rect 16390 7528 16396 7540
rect 2746 7500 16396 7528
rect 2148 7460 2176 7488
rect 2746 7460 2774 7500
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 19978 7528 19984 7540
rect 16592 7500 19984 7528
rect 2148 7432 2774 7460
rect 4798 7420 4804 7472
rect 4856 7460 4862 7472
rect 11054 7460 11060 7472
rect 4856 7432 11060 7460
rect 4856 7420 4862 7432
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 16592 7392 16620 7500
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 20162 7488 20168 7540
rect 20220 7488 20226 7540
rect 20346 7488 20352 7540
rect 20404 7528 20410 7540
rect 20625 7531 20683 7537
rect 20625 7528 20637 7531
rect 20404 7500 20637 7528
rect 20404 7488 20410 7500
rect 20625 7497 20637 7500
rect 20671 7497 20683 7531
rect 20625 7491 20683 7497
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 22370 7528 22376 7540
rect 20772 7500 22376 7528
rect 20772 7488 20778 7500
rect 22370 7488 22376 7500
rect 22428 7488 22434 7540
rect 22557 7531 22615 7537
rect 22557 7497 22569 7531
rect 22603 7528 22615 7531
rect 22646 7528 22652 7540
rect 22603 7500 22652 7528
rect 22603 7497 22615 7500
rect 22557 7491 22615 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 23109 7531 23167 7537
rect 23109 7497 23121 7531
rect 23155 7497 23167 7531
rect 23109 7491 23167 7497
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 17000 7432 20944 7460
rect 17000 7420 17006 7432
rect 1811 7364 16620 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 17184 7364 19748 7392
rect 17184 7352 17190 7364
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 16482 7324 16488 7336
rect 6972 7296 16488 7324
rect 6972 7284 6978 7296
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 19610 7284 19616 7336
rect 19668 7284 19674 7336
rect 19720 7324 19748 7364
rect 19794 7352 19800 7404
rect 19852 7352 19858 7404
rect 19978 7352 19984 7404
rect 20036 7352 20042 7404
rect 20254 7352 20260 7404
rect 20312 7392 20318 7404
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20312 7364 20545 7392
rect 20312 7352 20318 7364
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 20806 7352 20812 7404
rect 20864 7352 20870 7404
rect 20916 7392 20944 7432
rect 20916 7364 21128 7392
rect 19720 7296 20484 7324
rect 19628 7197 19656 7284
rect 19702 7216 19708 7268
rect 19760 7216 19766 7268
rect 19613 7191 19671 7197
rect 19613 7157 19625 7191
rect 19659 7157 19671 7191
rect 19720 7188 19748 7216
rect 20349 7191 20407 7197
rect 20349 7188 20361 7191
rect 19720 7160 20361 7188
rect 19613 7151 19671 7157
rect 20349 7157 20361 7160
rect 20395 7157 20407 7191
rect 20456 7188 20484 7296
rect 21100 7256 21128 7364
rect 22554 7352 22560 7404
rect 22612 7392 22618 7404
rect 22741 7395 22799 7401
rect 22741 7392 22753 7395
rect 22612 7364 22753 7392
rect 22612 7352 22618 7364
rect 22741 7361 22753 7364
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 21174 7284 21180 7336
rect 21232 7324 21238 7336
rect 23124 7324 23152 7491
rect 23290 7488 23296 7540
rect 23348 7488 23354 7540
rect 23382 7488 23388 7540
rect 23440 7528 23446 7540
rect 24673 7531 24731 7537
rect 24673 7528 24685 7531
rect 23440 7500 24685 7528
rect 23440 7488 23446 7500
rect 24673 7497 24685 7500
rect 24719 7497 24731 7531
rect 24673 7491 24731 7497
rect 24762 7488 24768 7540
rect 24820 7488 24826 7540
rect 24854 7488 24860 7540
rect 24912 7488 24918 7540
rect 25038 7488 25044 7540
rect 25096 7528 25102 7540
rect 28994 7528 29000 7540
rect 25096 7500 29000 7528
rect 25096 7488 25102 7500
rect 28994 7488 29000 7500
rect 29052 7488 29058 7540
rect 31386 7488 31392 7540
rect 31444 7488 31450 7540
rect 44542 7488 44548 7540
rect 44600 7528 44606 7540
rect 45097 7531 45155 7537
rect 45097 7528 45109 7531
rect 44600 7500 45109 7528
rect 44600 7488 44606 7500
rect 45097 7497 45109 7500
rect 45143 7497 45155 7531
rect 45097 7491 45155 7497
rect 45278 7488 45284 7540
rect 45336 7488 45342 7540
rect 45646 7488 45652 7540
rect 45704 7488 45710 7540
rect 46382 7488 46388 7540
rect 46440 7488 46446 7540
rect 23308 7460 23336 7488
rect 24780 7460 24808 7488
rect 23308 7432 24164 7460
rect 23293 7395 23351 7401
rect 23293 7361 23305 7395
rect 23339 7392 23351 7395
rect 23474 7392 23480 7404
rect 23339 7364 23480 7392
rect 23339 7361 23351 7364
rect 23293 7355 23351 7361
rect 23474 7352 23480 7364
rect 23532 7352 23538 7404
rect 23569 7395 23627 7401
rect 23569 7361 23581 7395
rect 23615 7392 23627 7395
rect 23658 7392 23664 7404
rect 23615 7364 23664 7392
rect 23615 7361 23627 7364
rect 23569 7355 23627 7361
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 23842 7352 23848 7404
rect 23900 7352 23906 7404
rect 21232 7296 23152 7324
rect 21232 7284 21238 7296
rect 23661 7259 23719 7265
rect 23661 7256 23673 7259
rect 21100 7228 23673 7256
rect 23661 7225 23673 7228
rect 23707 7225 23719 7259
rect 24136 7256 24164 7432
rect 24228 7432 24808 7460
rect 24872 7460 24900 7488
rect 31110 7460 31116 7472
rect 24872 7432 31116 7460
rect 24228 7401 24256 7432
rect 31110 7420 31116 7432
rect 31168 7420 31174 7472
rect 24213 7395 24271 7401
rect 24213 7361 24225 7395
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 24581 7395 24639 7401
rect 24581 7361 24593 7395
rect 24627 7361 24639 7395
rect 24581 7355 24639 7361
rect 24857 7395 24915 7401
rect 24857 7361 24869 7395
rect 24903 7392 24915 7395
rect 31404 7392 31432 7488
rect 44821 7463 44879 7469
rect 44821 7429 44833 7463
rect 44867 7460 44879 7463
rect 45296 7460 45324 7488
rect 44867 7432 45324 7460
rect 44867 7429 44879 7432
rect 44821 7423 44879 7429
rect 24903 7364 31432 7392
rect 24903 7361 24915 7364
rect 24857 7355 24915 7361
rect 24596 7324 24624 7355
rect 41598 7352 41604 7404
rect 41656 7392 41662 7404
rect 44453 7395 44511 7401
rect 44453 7392 44465 7395
rect 41656 7364 44465 7392
rect 41656 7352 41662 7364
rect 44453 7361 44465 7364
rect 44499 7361 44511 7395
rect 44453 7355 44511 7361
rect 45005 7395 45063 7401
rect 45005 7361 45017 7395
rect 45051 7361 45063 7395
rect 45005 7355 45063 7361
rect 29086 7324 29092 7336
rect 24596 7296 29092 7324
rect 29086 7284 29092 7296
rect 29144 7284 29150 7336
rect 36446 7284 36452 7336
rect 36504 7324 36510 7336
rect 45020 7324 45048 7355
rect 45554 7352 45560 7404
rect 45612 7352 45618 7404
rect 45646 7352 45652 7404
rect 45704 7392 45710 7404
rect 46109 7395 46167 7401
rect 46109 7392 46121 7395
rect 45704 7364 46121 7392
rect 45704 7352 45710 7364
rect 46109 7361 46121 7364
rect 46155 7361 46167 7395
rect 46109 7355 46167 7361
rect 36504 7296 45048 7324
rect 36504 7284 36510 7296
rect 36906 7256 36912 7268
rect 24136 7228 36912 7256
rect 23661 7219 23719 7225
rect 36906 7216 36912 7228
rect 36964 7216 36970 7268
rect 22738 7188 22744 7200
rect 20456 7160 22744 7188
rect 20349 7151 20407 7157
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 23382 7148 23388 7200
rect 23440 7148 23446 7200
rect 24026 7148 24032 7200
rect 24084 7148 24090 7200
rect 24397 7191 24455 7197
rect 24397 7157 24409 7191
rect 24443 7188 24455 7191
rect 24670 7188 24676 7200
rect 24443 7160 24676 7188
rect 24443 7157 24455 7160
rect 24397 7151 24455 7157
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 1104 7098 46828 7120
rect 1104 7046 6665 7098
rect 6717 7046 6729 7098
rect 6781 7046 6793 7098
rect 6845 7046 6857 7098
rect 6909 7046 6921 7098
rect 6973 7046 18095 7098
rect 18147 7046 18159 7098
rect 18211 7046 18223 7098
rect 18275 7046 18287 7098
rect 18339 7046 18351 7098
rect 18403 7046 29525 7098
rect 29577 7046 29589 7098
rect 29641 7046 29653 7098
rect 29705 7046 29717 7098
rect 29769 7046 29781 7098
rect 29833 7046 40955 7098
rect 41007 7046 41019 7098
rect 41071 7046 41083 7098
rect 41135 7046 41147 7098
rect 41199 7046 41211 7098
rect 41263 7046 46828 7098
rect 1104 7024 46828 7046
rect 15746 6944 15752 6996
rect 15804 6944 15810 6996
rect 17034 6944 17040 6996
rect 17092 6984 17098 6996
rect 21174 6984 21180 6996
rect 17092 6956 21180 6984
rect 17092 6944 17098 6956
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 21376 6956 23428 6984
rect 15764 6916 15792 6944
rect 21376 6916 21404 6956
rect 23400 6928 23428 6956
rect 23474 6944 23480 6996
rect 23532 6984 23538 6996
rect 28902 6984 28908 6996
rect 23532 6956 28908 6984
rect 23532 6944 23538 6956
rect 28902 6944 28908 6956
rect 28960 6944 28966 6996
rect 46014 6944 46020 6996
rect 46072 6984 46078 6996
rect 46201 6987 46259 6993
rect 46201 6984 46213 6987
rect 46072 6956 46213 6984
rect 46072 6944 46078 6956
rect 46201 6953 46213 6956
rect 46247 6953 46259 6987
rect 46201 6947 46259 6953
rect 15764 6888 21404 6916
rect 23382 6876 23388 6928
rect 23440 6876 23446 6928
rect 23842 6876 23848 6928
rect 23900 6916 23906 6928
rect 28442 6916 28448 6928
rect 23900 6888 28448 6916
rect 23900 6876 23906 6888
rect 28442 6876 28448 6888
rect 28500 6876 28506 6928
rect 15286 6808 15292 6860
rect 15344 6848 15350 6860
rect 22922 6848 22928 6860
rect 15344 6820 22928 6848
rect 15344 6808 15350 6820
rect 22922 6808 22928 6820
rect 22980 6808 22986 6860
rect 44910 6808 44916 6860
rect 44968 6848 44974 6860
rect 45833 6851 45891 6857
rect 45833 6848 45845 6851
rect 44968 6820 45845 6848
rect 44968 6808 44974 6820
rect 45833 6817 45845 6820
rect 45879 6817 45891 6851
rect 45833 6811 45891 6817
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 23198 6780 23204 6792
rect 16172 6752 23204 6780
rect 16172 6740 16178 6752
rect 23198 6740 23204 6752
rect 23256 6740 23262 6792
rect 44358 6740 44364 6792
rect 44416 6780 44422 6792
rect 46109 6783 46167 6789
rect 46109 6780 46121 6783
rect 44416 6752 46121 6780
rect 44416 6740 44422 6752
rect 46109 6749 46121 6752
rect 46155 6749 46167 6783
rect 46109 6743 46167 6749
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 22646 6712 22652 6724
rect 16540 6684 22652 6712
rect 16540 6672 16546 6684
rect 22646 6672 22652 6684
rect 22704 6672 22710 6724
rect 42794 6672 42800 6724
rect 42852 6712 42858 6724
rect 45557 6715 45615 6721
rect 45557 6712 45569 6715
rect 42852 6684 45569 6712
rect 42852 6672 42858 6684
rect 45557 6681 45569 6684
rect 45603 6681 45615 6715
rect 45557 6675 45615 6681
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 24026 6644 24032 6656
rect 9732 6616 24032 6644
rect 9732 6604 9738 6616
rect 24026 6604 24032 6616
rect 24084 6604 24090 6656
rect 1104 6554 46984 6576
rect 1104 6502 12380 6554
rect 12432 6502 12444 6554
rect 12496 6502 12508 6554
rect 12560 6502 12572 6554
rect 12624 6502 12636 6554
rect 12688 6502 23810 6554
rect 23862 6502 23874 6554
rect 23926 6502 23938 6554
rect 23990 6502 24002 6554
rect 24054 6502 24066 6554
rect 24118 6502 35240 6554
rect 35292 6502 35304 6554
rect 35356 6502 35368 6554
rect 35420 6502 35432 6554
rect 35484 6502 35496 6554
rect 35548 6502 46670 6554
rect 46722 6502 46734 6554
rect 46786 6502 46798 6554
rect 46850 6502 46862 6554
rect 46914 6502 46926 6554
rect 46978 6502 46984 6554
rect 1104 6480 46984 6502
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 25130 6440 25136 6452
rect 4396 6412 25136 6440
rect 4396 6400 4402 6412
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 25958 6372 25964 6384
rect 6512 6344 25964 6372
rect 6512 6332 6518 6344
rect 25958 6332 25964 6344
rect 26016 6332 26022 6384
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 24578 6304 24584 6316
rect 8352 6276 24584 6304
rect 8352 6264 8358 6276
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 20714 6236 20720 6248
rect 11112 6208 20720 6236
rect 11112 6196 11118 6208
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 24762 6128 24768 6180
rect 24820 6168 24826 6180
rect 34514 6168 34520 6180
rect 24820 6140 34520 6168
rect 24820 6128 24826 6140
rect 34514 6128 34520 6140
rect 34572 6128 34578 6180
rect 1104 6010 46828 6032
rect 1104 5958 6665 6010
rect 6717 5958 6729 6010
rect 6781 5958 6793 6010
rect 6845 5958 6857 6010
rect 6909 5958 6921 6010
rect 6973 5958 18095 6010
rect 18147 5958 18159 6010
rect 18211 5958 18223 6010
rect 18275 5958 18287 6010
rect 18339 5958 18351 6010
rect 18403 5958 29525 6010
rect 29577 5958 29589 6010
rect 29641 5958 29653 6010
rect 29705 5958 29717 6010
rect 29769 5958 29781 6010
rect 29833 5958 40955 6010
rect 41007 5958 41019 6010
rect 41071 5958 41083 6010
rect 41135 5958 41147 6010
rect 41199 5958 41211 6010
rect 41263 5958 46828 6010
rect 1104 5936 46828 5958
rect 32122 5584 32128 5636
rect 32180 5624 32186 5636
rect 36630 5624 36636 5636
rect 32180 5596 36636 5624
rect 32180 5584 32186 5596
rect 36630 5584 36636 5596
rect 36688 5584 36694 5636
rect 1104 5466 46984 5488
rect 1104 5414 12380 5466
rect 12432 5414 12444 5466
rect 12496 5414 12508 5466
rect 12560 5414 12572 5466
rect 12624 5414 12636 5466
rect 12688 5414 23810 5466
rect 23862 5414 23874 5466
rect 23926 5414 23938 5466
rect 23990 5414 24002 5466
rect 24054 5414 24066 5466
rect 24118 5414 35240 5466
rect 35292 5414 35304 5466
rect 35356 5414 35368 5466
rect 35420 5414 35432 5466
rect 35484 5414 35496 5466
rect 35548 5414 46670 5466
rect 46722 5414 46734 5466
rect 46786 5414 46798 5466
rect 46850 5414 46862 5466
rect 46914 5414 46926 5466
rect 46978 5414 46984 5466
rect 1104 5392 46984 5414
rect 24670 4972 24676 5024
rect 24728 5012 24734 5024
rect 34606 5012 34612 5024
rect 24728 4984 34612 5012
rect 24728 4972 24734 4984
rect 34606 4972 34612 4984
rect 34664 4972 34670 5024
rect 1104 4922 46828 4944
rect 1104 4870 6665 4922
rect 6717 4870 6729 4922
rect 6781 4870 6793 4922
rect 6845 4870 6857 4922
rect 6909 4870 6921 4922
rect 6973 4870 18095 4922
rect 18147 4870 18159 4922
rect 18211 4870 18223 4922
rect 18275 4870 18287 4922
rect 18339 4870 18351 4922
rect 18403 4870 29525 4922
rect 29577 4870 29589 4922
rect 29641 4870 29653 4922
rect 29705 4870 29717 4922
rect 29769 4870 29781 4922
rect 29833 4870 40955 4922
rect 41007 4870 41019 4922
rect 41071 4870 41083 4922
rect 41135 4870 41147 4922
rect 41199 4870 41211 4922
rect 41263 4870 46828 4922
rect 1104 4848 46828 4870
rect 27706 4768 27712 4820
rect 27764 4808 27770 4820
rect 45094 4808 45100 4820
rect 27764 4780 45100 4808
rect 27764 4768 27770 4780
rect 45094 4768 45100 4780
rect 45152 4768 45158 4820
rect 1104 4378 46984 4400
rect 1104 4326 12380 4378
rect 12432 4326 12444 4378
rect 12496 4326 12508 4378
rect 12560 4326 12572 4378
rect 12624 4326 12636 4378
rect 12688 4326 23810 4378
rect 23862 4326 23874 4378
rect 23926 4326 23938 4378
rect 23990 4326 24002 4378
rect 24054 4326 24066 4378
rect 24118 4326 35240 4378
rect 35292 4326 35304 4378
rect 35356 4326 35368 4378
rect 35420 4326 35432 4378
rect 35484 4326 35496 4378
rect 35548 4326 46670 4378
rect 46722 4326 46734 4378
rect 46786 4326 46798 4378
rect 46850 4326 46862 4378
rect 46914 4326 46926 4378
rect 46978 4326 46984 4378
rect 1104 4304 46984 4326
rect 1104 3834 46828 3856
rect 1104 3782 6665 3834
rect 6717 3782 6729 3834
rect 6781 3782 6793 3834
rect 6845 3782 6857 3834
rect 6909 3782 6921 3834
rect 6973 3782 18095 3834
rect 18147 3782 18159 3834
rect 18211 3782 18223 3834
rect 18275 3782 18287 3834
rect 18339 3782 18351 3834
rect 18403 3782 29525 3834
rect 29577 3782 29589 3834
rect 29641 3782 29653 3834
rect 29705 3782 29717 3834
rect 29769 3782 29781 3834
rect 29833 3782 40955 3834
rect 41007 3782 41019 3834
rect 41071 3782 41083 3834
rect 41135 3782 41147 3834
rect 41199 3782 41211 3834
rect 41263 3782 46828 3834
rect 1104 3760 46828 3782
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 33686 3652 33692 3664
rect 24268 3624 33692 3652
rect 24268 3612 24274 3624
rect 33686 3612 33692 3624
rect 33744 3612 33750 3664
rect 23658 3544 23664 3596
rect 23716 3584 23722 3596
rect 36078 3584 36084 3596
rect 23716 3556 36084 3584
rect 23716 3544 23722 3556
rect 36078 3544 36084 3556
rect 36136 3544 36142 3596
rect 29914 3476 29920 3528
rect 29972 3516 29978 3528
rect 43990 3516 43996 3528
rect 29972 3488 43996 3516
rect 29972 3476 29978 3488
rect 43990 3476 43996 3488
rect 44048 3476 44054 3528
rect 25682 3408 25688 3460
rect 25740 3448 25746 3460
rect 39942 3448 39948 3460
rect 25740 3420 39948 3448
rect 25740 3408 25746 3420
rect 39942 3408 39948 3420
rect 40000 3408 40006 3460
rect 1104 3290 46984 3312
rect 1104 3238 12380 3290
rect 12432 3238 12444 3290
rect 12496 3238 12508 3290
rect 12560 3238 12572 3290
rect 12624 3238 12636 3290
rect 12688 3238 23810 3290
rect 23862 3238 23874 3290
rect 23926 3238 23938 3290
rect 23990 3238 24002 3290
rect 24054 3238 24066 3290
rect 24118 3238 35240 3290
rect 35292 3238 35304 3290
rect 35356 3238 35368 3290
rect 35420 3238 35432 3290
rect 35484 3238 35496 3290
rect 35548 3238 46670 3290
rect 46722 3238 46734 3290
rect 46786 3238 46798 3290
rect 46850 3238 46862 3290
rect 46914 3238 46926 3290
rect 46978 3238 46984 3290
rect 1104 3216 46984 3238
rect 1104 2746 46828 2768
rect 1104 2694 6665 2746
rect 6717 2694 6729 2746
rect 6781 2694 6793 2746
rect 6845 2694 6857 2746
rect 6909 2694 6921 2746
rect 6973 2694 18095 2746
rect 18147 2694 18159 2746
rect 18211 2694 18223 2746
rect 18275 2694 18287 2746
rect 18339 2694 18351 2746
rect 18403 2694 29525 2746
rect 29577 2694 29589 2746
rect 29641 2694 29653 2746
rect 29705 2694 29717 2746
rect 29769 2694 29781 2746
rect 29833 2694 40955 2746
rect 41007 2694 41019 2746
rect 41071 2694 41083 2746
rect 41135 2694 41147 2746
rect 41199 2694 41211 2746
rect 41263 2694 46828 2746
rect 1104 2672 46828 2694
rect 23658 2592 23664 2644
rect 23716 2592 23722 2644
rect 24210 2592 24216 2644
rect 24268 2592 24274 2644
rect 24762 2592 24768 2644
rect 24820 2592 24826 2644
rect 25593 2635 25651 2641
rect 25593 2601 25605 2635
rect 25639 2632 25651 2635
rect 27614 2632 27620 2644
rect 25639 2604 27620 2632
rect 25639 2601 25651 2604
rect 25593 2595 25651 2601
rect 27614 2592 27620 2604
rect 27672 2592 27678 2644
rect 27706 2592 27712 2644
rect 27764 2592 27770 2644
rect 29914 2592 29920 2644
rect 29972 2592 29978 2644
rect 32122 2592 32128 2644
rect 32180 2592 32186 2644
rect 34333 2635 34391 2641
rect 34333 2601 34345 2635
rect 34379 2632 34391 2635
rect 36446 2632 36452 2644
rect 34379 2604 36452 2632
rect 34379 2601 34391 2604
rect 34333 2595 34391 2601
rect 36446 2592 36452 2604
rect 36504 2592 36510 2644
rect 38841 2635 38899 2641
rect 38841 2601 38853 2635
rect 38887 2632 38899 2635
rect 41598 2632 41604 2644
rect 38887 2604 41604 2632
rect 38887 2601 38899 2604
rect 38841 2595 38899 2601
rect 41598 2592 41604 2604
rect 41656 2592 41662 2644
rect 42794 2592 42800 2644
rect 42852 2592 42858 2644
rect 43257 2635 43315 2641
rect 43257 2601 43269 2635
rect 43303 2632 43315 2635
rect 44358 2632 44364 2644
rect 43303 2604 44364 2632
rect 43303 2601 43315 2604
rect 43257 2595 43315 2601
rect 44358 2592 44364 2604
rect 44416 2592 44422 2644
rect 45189 2635 45247 2641
rect 45189 2601 45201 2635
rect 45235 2632 45247 2635
rect 45554 2632 45560 2644
rect 45235 2604 45560 2632
rect 45235 2601 45247 2604
rect 45189 2595 45247 2601
rect 45554 2592 45560 2604
rect 45612 2592 45618 2644
rect 45646 2592 45652 2644
rect 45704 2592 45710 2644
rect 45738 2592 45744 2644
rect 45796 2592 45802 2644
rect 23474 2524 23480 2576
rect 23532 2564 23538 2576
rect 25041 2567 25099 2573
rect 23532 2536 24900 2564
rect 23532 2524 23538 2536
rect 23385 2499 23443 2505
rect 23385 2465 23397 2499
rect 23431 2496 23443 2499
rect 24762 2496 24768 2508
rect 23431 2468 24768 2496
rect 23431 2465 23443 2468
rect 23385 2459 23443 2465
rect 24762 2456 24768 2468
rect 24820 2456 24826 2508
rect 24872 2496 24900 2536
rect 25041 2533 25053 2567
rect 25087 2564 25099 2567
rect 25317 2567 25375 2573
rect 25087 2536 25268 2564
rect 25087 2533 25099 2536
rect 25041 2527 25099 2533
rect 25240 2496 25268 2536
rect 25317 2533 25329 2567
rect 25363 2564 25375 2567
rect 36633 2567 36691 2573
rect 25363 2536 35940 2564
rect 25363 2533 25375 2536
rect 25317 2527 25375 2533
rect 35912 2496 35940 2536
rect 36633 2533 36645 2567
rect 36679 2564 36691 2567
rect 42812 2564 42840 2592
rect 36679 2536 42840 2564
rect 36679 2533 36691 2536
rect 36633 2527 36691 2533
rect 40034 2496 40040 2508
rect 24872 2468 24992 2496
rect 25240 2468 35756 2496
rect 35912 2468 40040 2496
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 22428 2400 23489 2428
rect 22428 2388 22434 2400
rect 23477 2397 23489 2400
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 23753 2431 23811 2437
rect 23753 2428 23765 2431
rect 23716 2400 23765 2428
rect 23716 2388 23722 2400
rect 23753 2397 23765 2400
rect 23799 2397 23811 2431
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23753 2391 23811 2397
rect 23860 2400 24041 2428
rect 21082 2320 21088 2372
rect 21140 2320 21146 2372
rect 23198 2320 23204 2372
rect 23256 2320 23262 2372
rect 23566 2320 23572 2372
rect 23624 2360 23630 2372
rect 23860 2360 23888 2400
rect 24029 2397 24041 2400
rect 24075 2397 24087 2431
rect 24029 2391 24087 2397
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 24854 2388 24860 2440
rect 24912 2388 24918 2440
rect 24964 2428 24992 2468
rect 25133 2431 25191 2437
rect 25133 2428 25145 2431
rect 24964 2400 25145 2428
rect 25133 2397 25145 2400
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 25406 2388 25412 2440
rect 25464 2388 25470 2440
rect 27522 2388 27528 2440
rect 27580 2388 27586 2440
rect 29730 2388 29736 2440
rect 29788 2388 29794 2440
rect 31386 2388 31392 2440
rect 31444 2428 31450 2440
rect 31941 2431 31999 2437
rect 31941 2428 31953 2431
rect 31444 2400 31953 2428
rect 31444 2388 31450 2400
rect 31941 2397 31953 2400
rect 31987 2397 31999 2431
rect 31941 2391 31999 2397
rect 34146 2388 34152 2440
rect 34204 2388 34210 2440
rect 35728 2360 35756 2468
rect 40034 2456 40040 2468
rect 40092 2456 40098 2508
rect 40218 2456 40224 2508
rect 40276 2456 40282 2508
rect 36446 2388 36452 2440
rect 36504 2388 36510 2440
rect 38654 2388 38660 2440
rect 38712 2388 38718 2440
rect 40236 2360 40264 2456
rect 43070 2388 43076 2440
rect 43128 2388 43134 2440
rect 45002 2388 45008 2440
rect 45060 2388 45066 2440
rect 45465 2431 45523 2437
rect 45465 2397 45477 2431
rect 45511 2397 45523 2431
rect 45465 2391 45523 2397
rect 23624 2332 23888 2360
rect 24872 2332 35664 2360
rect 35728 2332 40264 2360
rect 23624 2320 23630 2332
rect 21174 2252 21180 2304
rect 21232 2252 21238 2304
rect 23937 2295 23995 2301
rect 23937 2261 23949 2295
rect 23983 2292 23995 2295
rect 24872 2292 24900 2332
rect 23983 2264 24900 2292
rect 23983 2261 23995 2264
rect 23937 2255 23995 2261
rect 24946 2252 24952 2304
rect 25004 2292 25010 2304
rect 33870 2292 33876 2304
rect 25004 2264 33876 2292
rect 25004 2252 25010 2264
rect 33870 2252 33876 2264
rect 33928 2252 33934 2304
rect 35636 2292 35664 2332
rect 40586 2320 40592 2372
rect 40644 2320 40650 2372
rect 44726 2320 44732 2372
rect 44784 2360 44790 2372
rect 45480 2360 45508 2391
rect 45922 2388 45928 2440
rect 45980 2388 45986 2440
rect 44784 2332 45508 2360
rect 44784 2320 44790 2332
rect 40604 2292 40632 2320
rect 35636 2264 40632 2292
rect 1104 2202 46984 2224
rect 1104 2150 12380 2202
rect 12432 2150 12444 2202
rect 12496 2150 12508 2202
rect 12560 2150 12572 2202
rect 12624 2150 12636 2202
rect 12688 2150 23810 2202
rect 23862 2150 23874 2202
rect 23926 2150 23938 2202
rect 23990 2150 24002 2202
rect 24054 2150 24066 2202
rect 24118 2150 35240 2202
rect 35292 2150 35304 2202
rect 35356 2150 35368 2202
rect 35420 2150 35432 2202
rect 35484 2150 35496 2202
rect 35548 2150 46670 2202
rect 46722 2150 46734 2202
rect 46786 2150 46798 2202
rect 46850 2150 46862 2202
rect 46914 2150 46926 2202
rect 46978 2150 46984 2202
rect 1104 2128 46984 2150
rect 20257 2091 20315 2097
rect 20257 2057 20269 2091
rect 20303 2088 20315 2091
rect 21082 2088 21088 2100
rect 20303 2060 21088 2088
rect 20303 2057 20315 2060
rect 20257 2051 20315 2057
rect 21082 2048 21088 2060
rect 21140 2048 21146 2100
rect 21174 2048 21180 2100
rect 21232 2048 21238 2100
rect 22370 2048 22376 2100
rect 22428 2048 22434 2100
rect 22649 2091 22707 2097
rect 22649 2057 22661 2091
rect 22695 2088 22707 2091
rect 23198 2088 23204 2100
rect 22695 2060 23204 2088
rect 22695 2057 22707 2060
rect 22649 2051 22707 2057
rect 23198 2048 23204 2060
rect 23256 2048 23262 2100
rect 23385 2091 23443 2097
rect 23385 2057 23397 2091
rect 23431 2088 23443 2091
rect 23474 2088 23480 2100
rect 23431 2060 23480 2088
rect 23431 2057 23443 2060
rect 23385 2051 23443 2057
rect 23474 2048 23480 2060
rect 23532 2048 23538 2100
rect 23937 2091 23995 2097
rect 23937 2057 23949 2091
rect 23983 2088 23995 2091
rect 24578 2088 24584 2100
rect 23983 2060 24584 2088
rect 23983 2057 23995 2060
rect 23937 2051 23995 2057
rect 24578 2048 24584 2060
rect 24636 2048 24642 2100
rect 24673 2091 24731 2097
rect 24673 2057 24685 2091
rect 24719 2088 24731 2091
rect 25406 2088 25412 2100
rect 24719 2060 25412 2088
rect 24719 2057 24731 2060
rect 24673 2051 24731 2057
rect 25406 2048 25412 2060
rect 25464 2048 25470 2100
rect 27157 2091 27215 2097
rect 27157 2057 27169 2091
rect 27203 2088 27215 2091
rect 27522 2088 27528 2100
rect 27203 2060 27528 2088
rect 27203 2057 27215 2060
rect 27157 2051 27215 2057
rect 27522 2048 27528 2060
rect 27580 2048 27586 2100
rect 29273 2091 29331 2097
rect 29273 2057 29285 2091
rect 29319 2088 29331 2091
rect 29730 2088 29736 2100
rect 29319 2060 29736 2088
rect 29319 2057 29331 2060
rect 29273 2051 29331 2057
rect 29730 2048 29736 2060
rect 29788 2048 29794 2100
rect 31386 2048 31392 2100
rect 31444 2048 31450 2100
rect 33689 2091 33747 2097
rect 33689 2057 33701 2091
rect 33735 2088 33747 2091
rect 34146 2088 34152 2100
rect 33735 2060 34152 2088
rect 33735 2057 33747 2060
rect 33689 2051 33747 2057
rect 34146 2048 34152 2060
rect 34204 2048 34210 2100
rect 35713 2091 35771 2097
rect 35713 2057 35725 2091
rect 35759 2088 35771 2091
rect 36446 2088 36452 2100
rect 35759 2060 36452 2088
rect 35759 2057 35771 2060
rect 35713 2051 35771 2057
rect 36446 2048 36452 2060
rect 36504 2048 36510 2100
rect 37921 2091 37979 2097
rect 37921 2057 37933 2091
rect 37967 2088 37979 2091
rect 38654 2088 38660 2100
rect 37967 2060 38660 2088
rect 37967 2057 37979 2060
rect 37921 2051 37979 2057
rect 38654 2048 38660 2060
rect 38712 2048 38718 2100
rect 42613 2091 42671 2097
rect 42613 2057 42625 2091
rect 42659 2088 42671 2091
rect 43070 2088 43076 2100
rect 42659 2060 43076 2088
rect 42659 2057 42671 2060
rect 42613 2051 42671 2057
rect 43070 2048 43076 2060
rect 43128 2048 43134 2100
rect 43254 2048 43260 2100
rect 43312 2048 43318 2100
rect 44269 2091 44327 2097
rect 44269 2057 44281 2091
rect 44315 2088 44327 2091
rect 45002 2088 45008 2100
rect 44315 2060 45008 2088
rect 44315 2057 44327 2060
rect 44269 2051 44327 2057
rect 45002 2048 45008 2060
rect 45060 2048 45066 2100
rect 45833 2091 45891 2097
rect 45833 2057 45845 2091
rect 45879 2088 45891 2091
rect 45922 2088 45928 2100
rect 45879 2060 45928 2088
rect 45879 2057 45891 2060
rect 45833 2051 45891 2057
rect 45922 2048 45928 2060
rect 45980 2048 45986 2100
rect 21192 2020 21220 2048
rect 43272 2020 43300 2048
rect 21192 1992 43300 2020
rect 20070 1912 20076 1964
rect 20128 1912 20134 1964
rect 20898 1912 20904 1964
rect 20956 1952 20962 1964
rect 22189 1955 22247 1961
rect 22189 1952 22201 1955
rect 20956 1924 22201 1952
rect 20956 1912 20962 1924
rect 22189 1921 22201 1924
rect 22235 1921 22247 1955
rect 22189 1915 22247 1921
rect 22462 1912 22468 1964
rect 22520 1912 22526 1964
rect 22922 1912 22928 1964
rect 22980 1912 22986 1964
rect 23201 1955 23259 1961
rect 23201 1921 23213 1955
rect 23247 1921 23259 1955
rect 23201 1915 23259 1921
rect 19886 1844 19892 1896
rect 19944 1884 19950 1896
rect 23216 1884 23244 1915
rect 23474 1912 23480 1964
rect 23532 1912 23538 1964
rect 23753 1955 23811 1961
rect 23753 1921 23765 1955
rect 23799 1921 23811 1955
rect 23753 1915 23811 1921
rect 19944 1856 23244 1884
rect 19944 1844 19950 1856
rect 23290 1844 23296 1896
rect 23348 1884 23354 1896
rect 23768 1884 23796 1915
rect 24026 1912 24032 1964
rect 24084 1912 24090 1964
rect 24486 1912 24492 1964
rect 24544 1912 24550 1964
rect 24762 1912 24768 1964
rect 24820 1912 24826 1964
rect 24854 1912 24860 1964
rect 24912 1912 24918 1964
rect 26970 1912 26976 1964
rect 27028 1912 27034 1964
rect 29086 1912 29092 1964
rect 29144 1912 29150 1964
rect 31202 1912 31208 1964
rect 31260 1912 31266 1964
rect 33502 1912 33508 1964
rect 33560 1912 33566 1964
rect 35526 1912 35532 1964
rect 35584 1912 35590 1964
rect 37734 1912 37740 1964
rect 37792 1912 37798 1964
rect 42426 1912 42432 1964
rect 42484 1912 42490 1964
rect 44082 1912 44088 1964
rect 44140 1912 44146 1964
rect 44542 1912 44548 1964
rect 44600 1912 44606 1964
rect 45646 1912 45652 1964
rect 45704 1912 45710 1964
rect 23348 1856 23796 1884
rect 23348 1844 23354 1856
rect 23109 1819 23167 1825
rect 23109 1785 23121 1819
rect 23155 1816 23167 1819
rect 23750 1816 23756 1828
rect 23155 1788 23756 1816
rect 23155 1785 23167 1788
rect 23109 1779 23167 1785
rect 23750 1776 23756 1788
rect 23808 1776 23814 1828
rect 24872 1816 24900 1912
rect 24136 1788 24900 1816
rect 23661 1751 23719 1757
rect 23661 1717 23673 1751
rect 23707 1748 23719 1751
rect 24136 1748 24164 1788
rect 25682 1776 25688 1828
rect 25740 1776 25746 1828
rect 44726 1776 44732 1828
rect 44784 1776 44790 1828
rect 23707 1720 24164 1748
rect 24213 1751 24271 1757
rect 23707 1717 23719 1720
rect 23661 1711 23719 1717
rect 24213 1717 24225 1751
rect 24259 1748 24271 1751
rect 24670 1748 24676 1760
rect 24259 1720 24676 1748
rect 24259 1717 24271 1720
rect 24213 1711 24271 1717
rect 24670 1708 24676 1720
rect 24728 1708 24734 1760
rect 24949 1751 25007 1757
rect 24949 1717 24961 1751
rect 24995 1748 25007 1751
rect 25700 1748 25728 1776
rect 24995 1720 25728 1748
rect 24995 1717 25007 1720
rect 24949 1711 25007 1717
rect 27614 1708 27620 1760
rect 27672 1748 27678 1760
rect 36814 1748 36820 1760
rect 27672 1720 36820 1748
rect 27672 1708 27678 1720
rect 36814 1708 36820 1720
rect 36872 1708 36878 1760
rect 1104 1658 46828 1680
rect 1104 1606 6665 1658
rect 6717 1606 6729 1658
rect 6781 1606 6793 1658
rect 6845 1606 6857 1658
rect 6909 1606 6921 1658
rect 6973 1606 18095 1658
rect 18147 1606 18159 1658
rect 18211 1606 18223 1658
rect 18275 1606 18287 1658
rect 18339 1606 18351 1658
rect 18403 1606 29525 1658
rect 29577 1606 29589 1658
rect 29641 1606 29653 1658
rect 29705 1606 29717 1658
rect 29769 1606 29781 1658
rect 29833 1606 40955 1658
rect 41007 1606 41019 1658
rect 41071 1606 41083 1658
rect 41135 1606 41147 1658
rect 41199 1606 41211 1658
rect 41263 1606 46828 1658
rect 1104 1584 46828 1606
rect 19797 1547 19855 1553
rect 19797 1513 19809 1547
rect 19843 1544 19855 1547
rect 20070 1544 20076 1556
rect 19843 1516 20076 1544
rect 19843 1513 19855 1516
rect 19797 1507 19855 1513
rect 20070 1504 20076 1516
rect 20128 1504 20134 1556
rect 22005 1547 22063 1553
rect 22005 1513 22017 1547
rect 22051 1544 22063 1547
rect 22462 1544 22468 1556
rect 22051 1516 22468 1544
rect 22051 1513 22063 1516
rect 22005 1507 22063 1513
rect 22462 1504 22468 1516
rect 22520 1504 22526 1556
rect 23566 1504 23572 1556
rect 23624 1544 23630 1556
rect 23661 1547 23719 1553
rect 23661 1544 23673 1547
rect 23624 1516 23673 1544
rect 23624 1504 23630 1516
rect 23661 1513 23673 1516
rect 23707 1513 23719 1547
rect 23661 1507 23719 1513
rect 24026 1504 24032 1556
rect 24084 1504 24090 1556
rect 24213 1547 24271 1553
rect 24213 1513 24225 1547
rect 24259 1544 24271 1547
rect 24486 1544 24492 1556
rect 24259 1516 24492 1544
rect 24259 1513 24271 1516
rect 24213 1507 24271 1513
rect 24486 1504 24492 1516
rect 24544 1504 24550 1556
rect 26421 1547 26479 1553
rect 26421 1513 26433 1547
rect 26467 1544 26479 1547
rect 26970 1544 26976 1556
rect 26467 1516 26976 1544
rect 26467 1513 26479 1516
rect 26421 1507 26479 1513
rect 26970 1504 26976 1516
rect 27028 1504 27034 1556
rect 28629 1547 28687 1553
rect 28629 1513 28641 1547
rect 28675 1544 28687 1547
rect 29086 1544 29092 1556
rect 28675 1516 29092 1544
rect 28675 1513 28687 1516
rect 28629 1507 28687 1513
rect 29086 1504 29092 1516
rect 29144 1504 29150 1556
rect 30837 1547 30895 1553
rect 30837 1513 30849 1547
rect 30883 1544 30895 1547
rect 31202 1544 31208 1556
rect 30883 1516 31208 1544
rect 30883 1513 30895 1516
rect 30837 1507 30895 1513
rect 31202 1504 31208 1516
rect 31260 1504 31266 1556
rect 33045 1547 33103 1553
rect 33045 1513 33057 1547
rect 33091 1544 33103 1547
rect 33502 1544 33508 1556
rect 33091 1516 33508 1544
rect 33091 1513 33103 1516
rect 33045 1507 33103 1513
rect 33502 1504 33508 1516
rect 33560 1504 33566 1556
rect 35253 1547 35311 1553
rect 35253 1513 35265 1547
rect 35299 1544 35311 1547
rect 35526 1544 35532 1556
rect 35299 1516 35532 1544
rect 35299 1513 35311 1516
rect 35253 1507 35311 1513
rect 35526 1504 35532 1516
rect 35584 1504 35590 1556
rect 37461 1547 37519 1553
rect 37461 1513 37473 1547
rect 37507 1544 37519 1547
rect 37734 1544 37740 1556
rect 37507 1516 37740 1544
rect 37507 1513 37519 1516
rect 37461 1507 37519 1513
rect 37734 1504 37740 1516
rect 37792 1504 37798 1556
rect 41877 1547 41935 1553
rect 41877 1513 41889 1547
rect 41923 1544 41935 1547
rect 42426 1544 42432 1556
rect 41923 1516 42432 1544
rect 41923 1513 41935 1516
rect 41877 1507 41935 1513
rect 42426 1504 42432 1516
rect 42484 1504 42490 1556
rect 44085 1547 44143 1553
rect 44085 1513 44097 1547
rect 44131 1544 44143 1547
rect 44542 1544 44548 1556
rect 44131 1516 44548 1544
rect 44131 1513 44143 1516
rect 44085 1507 44143 1513
rect 44542 1504 44548 1516
rect 44600 1504 44606 1556
rect 45646 1504 45652 1556
rect 45704 1544 45710 1556
rect 46109 1547 46167 1553
rect 46109 1544 46121 1547
rect 45704 1516 46121 1544
rect 45704 1504 45710 1516
rect 46109 1513 46121 1516
rect 46155 1513 46167 1547
rect 46109 1507 46167 1513
rect 15378 1436 15384 1488
rect 15436 1436 15442 1488
rect 23385 1479 23443 1485
rect 23385 1445 23397 1479
rect 23431 1476 23443 1479
rect 24044 1476 24072 1504
rect 23431 1448 24072 1476
rect 23431 1445 23443 1448
rect 23385 1439 23443 1445
rect 1946 1300 1952 1352
rect 2004 1300 2010 1352
rect 4154 1300 4160 1352
rect 4212 1300 4218 1352
rect 6362 1300 6368 1352
rect 6420 1300 6426 1352
rect 8570 1300 8576 1352
rect 8628 1300 8634 1352
rect 10778 1300 10784 1352
rect 10836 1300 10842 1352
rect 12986 1300 12992 1352
rect 13044 1300 13050 1352
rect 15194 1300 15200 1352
rect 15252 1300 15258 1352
rect 17402 1300 17408 1352
rect 17460 1300 17466 1352
rect 19610 1300 19616 1352
rect 19668 1300 19674 1352
rect 19996 1312 21128 1340
rect 19996 1272 20024 1312
rect 4356 1244 20024 1272
rect 2130 1164 2136 1216
rect 2188 1164 2194 1216
rect 4356 1213 4384 1244
rect 20898 1232 20904 1284
rect 20956 1232 20962 1284
rect 4341 1207 4399 1213
rect 4341 1173 4353 1207
rect 4387 1173 4399 1207
rect 4341 1167 4399 1173
rect 6546 1164 6552 1216
rect 6604 1164 6610 1216
rect 8754 1164 8760 1216
rect 8812 1164 8818 1216
rect 10962 1164 10968 1216
rect 11020 1164 11026 1216
rect 13173 1207 13231 1213
rect 13173 1173 13185 1207
rect 13219 1204 13231 1207
rect 15470 1204 15476 1216
rect 13219 1176 15476 1204
rect 13219 1173 13231 1176
rect 13173 1167 13231 1173
rect 15470 1164 15476 1176
rect 15528 1164 15534 1216
rect 17589 1207 17647 1213
rect 17589 1173 17601 1207
rect 17635 1204 17647 1207
rect 20916 1204 20944 1232
rect 17635 1176 20944 1204
rect 21100 1204 21128 1312
rect 21818 1300 21824 1352
rect 21876 1300 21882 1352
rect 23198 1300 23204 1352
rect 23256 1300 23262 1352
rect 23477 1343 23535 1349
rect 23477 1309 23489 1343
rect 23523 1309 23535 1343
rect 23477 1303 23535 1309
rect 21174 1232 21180 1284
rect 21232 1272 21238 1284
rect 23492 1272 23520 1303
rect 24026 1300 24032 1352
rect 24084 1300 24090 1352
rect 26234 1300 26240 1352
rect 26292 1300 26298 1352
rect 28442 1300 28448 1352
rect 28500 1300 28506 1352
rect 30650 1300 30656 1352
rect 30708 1300 30714 1352
rect 32858 1300 32864 1352
rect 32916 1300 32922 1352
rect 35066 1300 35072 1352
rect 35124 1300 35130 1352
rect 37274 1300 37280 1352
rect 37332 1300 37338 1352
rect 39482 1300 39488 1352
rect 39540 1300 39546 1352
rect 41690 1300 41696 1352
rect 41748 1300 41754 1352
rect 43898 1300 43904 1352
rect 43956 1300 43962 1352
rect 46290 1300 46296 1352
rect 46348 1300 46354 1352
rect 21232 1244 23520 1272
rect 21232 1232 21238 1244
rect 23474 1204 23480 1216
rect 21100 1176 23480 1204
rect 17635 1173 17647 1176
rect 17589 1167 17647 1173
rect 23474 1164 23480 1176
rect 23532 1164 23538 1216
rect 39669 1207 39727 1213
rect 39669 1173 39681 1207
rect 39715 1204 39727 1207
rect 44082 1204 44088 1216
rect 39715 1176 44088 1204
rect 39715 1173 39727 1176
rect 39669 1167 39727 1173
rect 44082 1164 44088 1176
rect 44140 1164 44146 1216
rect 1104 1114 46984 1136
rect 1104 1062 12380 1114
rect 12432 1062 12444 1114
rect 12496 1062 12508 1114
rect 12560 1062 12572 1114
rect 12624 1062 12636 1114
rect 12688 1062 23810 1114
rect 23862 1062 23874 1114
rect 23926 1062 23938 1114
rect 23990 1062 24002 1114
rect 24054 1062 24066 1114
rect 24118 1062 35240 1114
rect 35292 1062 35304 1114
rect 35356 1062 35368 1114
rect 35420 1062 35432 1114
rect 35484 1062 35496 1114
rect 35548 1062 46670 1114
rect 46722 1062 46734 1114
rect 46786 1062 46798 1114
rect 46850 1062 46862 1114
rect 46914 1062 46926 1114
rect 46978 1062 46984 1114
rect 1104 1040 46984 1062
rect 2130 960 2136 1012
rect 2188 1000 2194 1012
rect 2188 972 6914 1000
rect 2188 960 2194 972
rect 6546 892 6552 944
rect 6604 892 6610 944
rect 6564 728 6592 892
rect 6886 796 6914 972
rect 8754 960 8760 1012
rect 8812 1000 8818 1012
rect 19886 1000 19892 1012
rect 8812 972 19892 1000
rect 8812 960 8818 972
rect 19886 960 19892 972
rect 19944 960 19950 1012
rect 21174 960 21180 1012
rect 21232 960 21238 1012
rect 23198 960 23204 1012
rect 23256 960 23262 1012
rect 15378 892 15384 944
rect 15436 892 15442 944
rect 15470 892 15476 944
rect 15528 932 15534 944
rect 21192 932 21220 960
rect 15528 904 21220 932
rect 15528 892 15534 904
rect 15396 864 15424 892
rect 23216 864 23244 960
rect 15396 836 23244 864
rect 24762 796 24768 808
rect 6886 768 24768 796
rect 24762 756 24768 768
rect 24820 756 24826 808
rect 6564 700 6914 728
rect 6886 660 6914 700
rect 10962 688 10968 740
rect 11020 728 11026 740
rect 23290 728 23296 740
rect 11020 700 23296 728
rect 11020 688 11026 700
rect 23290 688 23296 700
rect 23348 688 23354 740
rect 22922 660 22928 672
rect 6886 632 22928 660
rect 22922 620 22928 632
rect 22980 620 22986 672
<< via1 >>
rect 7196 9936 7248 9988
rect 16856 9936 16908 9988
rect 10140 9868 10192 9920
rect 21548 9936 21600 9988
rect 24032 9936 24084 9988
rect 35072 9936 35124 9988
rect 12716 9800 12768 9852
rect 16120 9800 16172 9852
rect 20720 9868 20772 9920
rect 20904 9868 20956 9920
rect 22284 9868 22336 9920
rect 11888 9664 11940 9716
rect 22192 9800 22244 9852
rect 28816 9868 28868 9920
rect 28908 9868 28960 9920
rect 17408 9732 17460 9784
rect 24400 9800 24452 9852
rect 17868 9664 17920 9716
rect 27068 9732 27120 9784
rect 22652 9664 22704 9716
rect 24216 9664 24268 9716
rect 6184 9596 6236 9648
rect 10048 9596 10100 9648
rect 17132 9528 17184 9580
rect 17776 9596 17828 9648
rect 19984 9596 20036 9648
rect 22192 9596 22244 9648
rect 24124 9596 24176 9648
rect 29276 9664 29328 9716
rect 34336 9664 34388 9716
rect 23480 9528 23532 9580
rect 23572 9528 23624 9580
rect 24400 9528 24452 9580
rect 18604 9460 18656 9512
rect 21824 9460 21876 9512
rect 22008 9460 22060 9512
rect 37648 9596 37700 9648
rect 24676 9528 24728 9580
rect 24768 9460 24820 9512
rect 28172 9528 28224 9580
rect 33232 9528 33284 9580
rect 7288 9188 7340 9240
rect 5356 9120 5408 9172
rect 12716 9392 12768 9444
rect 12808 9392 12860 9444
rect 17408 9392 17460 9444
rect 26516 9392 26568 9444
rect 33600 9460 33652 9512
rect 24860 9324 24912 9376
rect 27804 9324 27856 9376
rect 32588 9324 32640 9376
rect 33876 9324 33928 9376
rect 43812 9324 43864 9376
rect 4988 9052 5040 9104
rect 13636 9256 13688 9308
rect 22376 9256 22428 9308
rect 28356 9256 28408 9308
rect 34060 9256 34112 9308
rect 34612 9256 34664 9308
rect 42800 9256 42852 9308
rect 9128 9188 9180 9240
rect 21364 9188 21416 9240
rect 21456 9188 21508 9240
rect 22192 9188 22244 9240
rect 11980 9120 12032 9172
rect 12072 9120 12124 9172
rect 21640 9120 21692 9172
rect 10232 8984 10284 9036
rect 10508 8916 10560 8968
rect 12072 8916 12124 8968
rect 8484 8848 8536 8900
rect 13636 8984 13688 9036
rect 17224 9052 17276 9104
rect 20352 9052 20404 9104
rect 26884 9188 26936 9240
rect 28448 9188 28500 9240
rect 39120 9188 39172 9240
rect 27988 9120 28040 9172
rect 33968 9120 34020 9172
rect 34336 9120 34388 9172
rect 36452 9120 36504 9172
rect 21640 8984 21692 9036
rect 22468 9052 22520 9104
rect 25504 9052 25556 9104
rect 29092 9052 29144 9104
rect 32128 9052 32180 9104
rect 36636 9052 36688 9104
rect 45468 9052 45520 9104
rect 22744 8984 22796 9036
rect 24676 8984 24728 9036
rect 23112 8916 23164 8968
rect 36544 8984 36596 9036
rect 36820 8984 36872 9036
rect 45100 8984 45152 9036
rect 28356 8916 28408 8968
rect 37004 8916 37056 8968
rect 13360 8848 13412 8900
rect 13544 8848 13596 8900
rect 22008 8848 22060 8900
rect 22468 8848 22520 8900
rect 24860 8848 24912 8900
rect 1952 8780 2004 8832
rect 4712 8780 4764 8832
rect 9680 8780 9732 8832
rect 10600 8780 10652 8832
rect 23020 8780 23072 8832
rect 24124 8780 24176 8832
rect 27620 8780 27672 8832
rect 27804 8780 27856 8832
rect 36176 8848 36228 8900
rect 36268 8848 36320 8900
rect 43628 8848 43680 8900
rect 34520 8780 34572 8832
rect 40684 8780 40736 8832
rect 12380 8678 12432 8730
rect 12444 8678 12496 8730
rect 12508 8678 12560 8730
rect 12572 8678 12624 8730
rect 12636 8678 12688 8730
rect 23810 8678 23862 8730
rect 23874 8678 23926 8730
rect 23938 8678 23990 8730
rect 24002 8678 24054 8730
rect 24066 8678 24118 8730
rect 35240 8678 35292 8730
rect 35304 8678 35356 8730
rect 35368 8678 35420 8730
rect 35432 8678 35484 8730
rect 35496 8678 35548 8730
rect 46670 8678 46722 8730
rect 46734 8678 46786 8730
rect 46798 8678 46850 8730
rect 46862 8678 46914 8730
rect 46926 8678 46978 8730
rect 2228 8576 2280 8628
rect 2964 8576 3016 8628
rect 3332 8576 3384 8628
rect 3700 8576 3752 8628
rect 4436 8576 4488 8628
rect 4896 8576 4948 8628
rect 4988 8576 5040 8628
rect 5448 8576 5500 8628
rect 5908 8576 5960 8628
rect 6276 8576 6328 8628
rect 6736 8619 6788 8628
rect 6736 8585 6745 8619
rect 6745 8585 6779 8619
rect 6779 8585 6788 8619
rect 6736 8576 6788 8585
rect 7748 8576 7800 8628
rect 8208 8576 8260 8628
rect 8484 8576 8536 8628
rect 5356 8508 5408 8560
rect 8852 8576 8904 8628
rect 9496 8576 9548 8628
rect 10416 8576 10468 8628
rect 10968 8576 11020 8628
rect 11428 8576 11480 8628
rect 12164 8576 12216 8628
rect 12256 8619 12308 8628
rect 12256 8585 12265 8619
rect 12265 8585 12299 8619
rect 12299 8585 12308 8619
rect 12256 8576 12308 8585
rect 13268 8576 13320 8628
rect 14004 8576 14056 8628
rect 14924 8576 14976 8628
rect 15476 8576 15528 8628
rect 16212 8576 16264 8628
rect 16488 8576 16540 8628
rect 17316 8576 17368 8628
rect 17684 8576 17736 8628
rect 18052 8619 18104 8628
rect 18052 8585 18061 8619
rect 18061 8585 18095 8619
rect 18095 8585 18104 8619
rect 18052 8576 18104 8585
rect 18420 8576 18472 8628
rect 18788 8576 18840 8628
rect 19892 8576 19944 8628
rect 20352 8576 20404 8628
rect 20536 8576 20588 8628
rect 9588 8508 9640 8560
rect 10508 8508 10560 8560
rect 14832 8508 14884 8560
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 2596 8372 2648 8424
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 7196 8440 7248 8492
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7932 8372 7984 8424
rect 6460 8304 6512 8356
rect 7840 8304 7892 8356
rect 9128 8440 9180 8492
rect 10048 8440 10100 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 10600 8440 10652 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12808 8440 12860 8492
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 13544 8440 13596 8492
rect 14648 8440 14700 8492
rect 17132 8508 17184 8560
rect 19248 8551 19300 8560
rect 19248 8517 19257 8551
rect 19257 8517 19291 8551
rect 19291 8517 19300 8551
rect 19248 8508 19300 8517
rect 21456 8576 21508 8628
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 17040 8440 17092 8492
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 20168 8440 20220 8492
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 21732 8508 21784 8560
rect 21824 8440 21876 8492
rect 22284 8576 22336 8628
rect 22560 8576 22612 8628
rect 22652 8576 22704 8628
rect 23020 8576 23072 8628
rect 25780 8576 25832 8628
rect 30748 8576 30800 8628
rect 31116 8576 31168 8628
rect 32128 8619 32180 8628
rect 32128 8585 32137 8619
rect 32137 8585 32171 8619
rect 32171 8585 32180 8619
rect 32128 8576 32180 8585
rect 22560 8440 22612 8492
rect 23204 8508 23256 8560
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 23756 8508 23808 8560
rect 23848 8440 23900 8492
rect 24308 8508 24360 8560
rect 27344 8508 27396 8560
rect 30380 8508 30432 8560
rect 24400 8440 24452 8492
rect 19524 8372 19576 8424
rect 13452 8304 13504 8356
rect 14464 8304 14516 8356
rect 17224 8304 17276 8356
rect 19708 8304 19760 8356
rect 23756 8372 23808 8424
rect 24952 8483 25004 8492
rect 24952 8449 24961 8483
rect 24961 8449 24995 8483
rect 24995 8449 25004 8483
rect 24952 8440 25004 8449
rect 25320 8483 25372 8492
rect 25320 8449 25329 8483
rect 25329 8449 25363 8483
rect 25363 8449 25372 8483
rect 25320 8440 25372 8449
rect 25688 8483 25740 8492
rect 25688 8449 25697 8483
rect 25697 8449 25731 8483
rect 25731 8449 25740 8483
rect 25688 8440 25740 8449
rect 26056 8483 26108 8492
rect 26056 8449 26065 8483
rect 26065 8449 26099 8483
rect 26099 8449 26108 8483
rect 26056 8440 26108 8449
rect 26424 8483 26476 8492
rect 26424 8449 26433 8483
rect 26433 8449 26467 8483
rect 26467 8449 26476 8483
rect 26424 8440 26476 8449
rect 26792 8483 26844 8492
rect 26792 8449 26801 8483
rect 26801 8449 26835 8483
rect 26835 8449 26844 8483
rect 26792 8440 26844 8449
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 27528 8483 27580 8492
rect 27528 8449 27537 8483
rect 27537 8449 27571 8483
rect 27571 8449 27580 8483
rect 27528 8440 27580 8449
rect 27896 8483 27948 8492
rect 27896 8449 27905 8483
rect 27905 8449 27939 8483
rect 27939 8449 27948 8483
rect 27896 8440 27948 8449
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 28632 8483 28684 8492
rect 28632 8449 28641 8483
rect 28641 8449 28675 8483
rect 28675 8449 28684 8483
rect 28632 8440 28684 8449
rect 28724 8440 28776 8492
rect 29368 8483 29420 8492
rect 29368 8449 29377 8483
rect 29377 8449 29411 8483
rect 29411 8449 29420 8483
rect 29368 8440 29420 8449
rect 29736 8483 29788 8492
rect 29736 8449 29745 8483
rect 29745 8449 29779 8483
rect 29779 8449 29788 8483
rect 29736 8440 29788 8449
rect 30104 8483 30156 8492
rect 30104 8449 30113 8483
rect 30113 8449 30147 8483
rect 30147 8449 30156 8483
rect 30104 8440 30156 8449
rect 30196 8440 30248 8492
rect 31208 8483 31260 8492
rect 31208 8449 31217 8483
rect 31217 8449 31251 8483
rect 31251 8449 31260 8483
rect 31208 8440 31260 8449
rect 31576 8483 31628 8492
rect 31576 8449 31585 8483
rect 31585 8449 31619 8483
rect 31619 8449 31628 8483
rect 31576 8440 31628 8449
rect 31668 8440 31720 8492
rect 32312 8483 32364 8492
rect 32312 8449 32321 8483
rect 32321 8449 32355 8483
rect 32355 8449 32364 8483
rect 32312 8440 32364 8449
rect 32588 8576 32640 8628
rect 33232 8619 33284 8628
rect 33232 8585 33241 8619
rect 33241 8585 33275 8619
rect 33275 8585 33284 8619
rect 33232 8576 33284 8585
rect 33600 8619 33652 8628
rect 33600 8585 33609 8619
rect 33609 8585 33643 8619
rect 33643 8585 33652 8619
rect 33600 8576 33652 8585
rect 33968 8619 34020 8628
rect 33968 8585 33977 8619
rect 33977 8585 34011 8619
rect 34011 8585 34020 8619
rect 33968 8576 34020 8585
rect 34060 8576 34112 8628
rect 35072 8576 35124 8628
rect 36176 8619 36228 8628
rect 36176 8585 36185 8619
rect 36185 8585 36219 8619
rect 36219 8585 36228 8619
rect 36176 8576 36228 8585
rect 36544 8619 36596 8628
rect 36544 8585 36553 8619
rect 36553 8585 36587 8619
rect 36587 8585 36596 8619
rect 36544 8576 36596 8585
rect 36912 8576 36964 8628
rect 39120 8619 39172 8628
rect 39120 8585 39129 8619
rect 39129 8585 39163 8619
rect 39163 8585 39172 8619
rect 39120 8576 39172 8585
rect 39396 8576 39448 8628
rect 39764 8508 39816 8560
rect 40684 8576 40736 8628
rect 40868 8576 40920 8628
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 32680 8440 32732 8449
rect 33048 8483 33100 8492
rect 33048 8449 33057 8483
rect 33057 8449 33091 8483
rect 33091 8449 33100 8483
rect 33048 8440 33100 8449
rect 33416 8483 33468 8492
rect 33416 8449 33425 8483
rect 33425 8449 33459 8483
rect 33459 8449 33468 8483
rect 33416 8440 33468 8449
rect 33784 8483 33836 8492
rect 33784 8449 33793 8483
rect 33793 8449 33827 8483
rect 33827 8449 33836 8483
rect 33784 8440 33836 8449
rect 34152 8483 34204 8492
rect 34152 8449 34161 8483
rect 34161 8449 34195 8483
rect 34195 8449 34204 8483
rect 34152 8440 34204 8449
rect 34244 8440 34296 8492
rect 34888 8483 34940 8492
rect 34888 8449 34897 8483
rect 34897 8449 34931 8483
rect 34931 8449 34940 8483
rect 34888 8440 34940 8449
rect 34980 8440 35032 8492
rect 35624 8483 35676 8492
rect 35624 8449 35633 8483
rect 35633 8449 35667 8483
rect 35667 8449 35676 8483
rect 35624 8440 35676 8449
rect 35716 8440 35768 8492
rect 36360 8483 36412 8492
rect 36360 8449 36369 8483
rect 36369 8449 36403 8483
rect 36403 8449 36412 8483
rect 36360 8440 36412 8449
rect 36728 8483 36780 8492
rect 36728 8449 36737 8483
rect 36737 8449 36771 8483
rect 36771 8449 36780 8483
rect 36728 8440 36780 8449
rect 37096 8483 37148 8492
rect 37096 8449 37105 8483
rect 37105 8449 37139 8483
rect 37139 8449 37148 8483
rect 37096 8440 37148 8449
rect 37188 8440 37240 8492
rect 37832 8483 37884 8492
rect 37832 8449 37841 8483
rect 37841 8449 37875 8483
rect 37875 8449 37884 8483
rect 37832 8440 37884 8449
rect 38200 8483 38252 8492
rect 38200 8449 38209 8483
rect 38209 8449 38243 8483
rect 38243 8449 38252 8483
rect 38200 8440 38252 8449
rect 38568 8483 38620 8492
rect 38568 8449 38577 8483
rect 38577 8449 38611 8483
rect 38611 8449 38620 8483
rect 38568 8440 38620 8449
rect 38936 8483 38988 8492
rect 38936 8449 38945 8483
rect 38945 8449 38979 8483
rect 38979 8449 38988 8483
rect 38936 8440 38988 8449
rect 39304 8483 39356 8492
rect 39304 8449 39313 8483
rect 39313 8449 39347 8483
rect 39347 8449 39356 8483
rect 39304 8440 39356 8449
rect 39948 8483 40000 8492
rect 39948 8449 39957 8483
rect 39957 8449 39991 8483
rect 39991 8449 40000 8483
rect 39948 8440 40000 8449
rect 40224 8440 40276 8492
rect 40592 8440 40644 8492
rect 41236 8508 41288 8560
rect 42708 8576 42760 8628
rect 44456 8576 44508 8628
rect 42800 8508 42852 8560
rect 43352 8508 43404 8560
rect 22284 8304 22336 8356
rect 26148 8304 26200 8356
rect 27436 8304 27488 8356
rect 20720 8236 20772 8288
rect 21180 8279 21232 8288
rect 21180 8245 21189 8279
rect 21189 8245 21223 8279
rect 21223 8245 21232 8279
rect 21180 8236 21232 8245
rect 21456 8279 21508 8288
rect 21456 8245 21465 8279
rect 21465 8245 21499 8279
rect 21499 8245 21508 8279
rect 21456 8236 21508 8245
rect 21824 8279 21876 8288
rect 21824 8245 21833 8279
rect 21833 8245 21867 8279
rect 21867 8245 21876 8279
rect 21824 8236 21876 8245
rect 22008 8236 22060 8288
rect 22560 8279 22612 8288
rect 22560 8245 22569 8279
rect 22569 8245 22603 8279
rect 22603 8245 22612 8279
rect 22560 8236 22612 8245
rect 22652 8279 22704 8288
rect 22652 8245 22661 8279
rect 22661 8245 22695 8279
rect 22695 8245 22704 8279
rect 22652 8236 22704 8245
rect 22744 8236 22796 8288
rect 23572 8236 23624 8288
rect 24768 8279 24820 8288
rect 24768 8245 24777 8279
rect 24777 8245 24811 8279
rect 24811 8245 24820 8279
rect 24768 8236 24820 8245
rect 25136 8279 25188 8288
rect 25136 8245 25145 8279
rect 25145 8245 25179 8279
rect 25179 8245 25188 8279
rect 25136 8236 25188 8245
rect 25228 8236 25280 8288
rect 25872 8279 25924 8288
rect 25872 8245 25881 8279
rect 25881 8245 25915 8279
rect 25915 8245 25924 8279
rect 25872 8236 25924 8245
rect 26608 8279 26660 8288
rect 26608 8245 26617 8279
rect 26617 8245 26651 8279
rect 26651 8245 26660 8279
rect 26608 8236 26660 8245
rect 26792 8236 26844 8288
rect 27160 8236 27212 8288
rect 27528 8236 27580 8288
rect 29000 8304 29052 8356
rect 33692 8372 33744 8424
rect 43628 8483 43680 8492
rect 43628 8449 43637 8483
rect 43637 8449 43671 8483
rect 43671 8449 43680 8483
rect 43628 8440 43680 8449
rect 43812 8440 43864 8492
rect 45100 8483 45152 8492
rect 45100 8449 45109 8483
rect 45109 8449 45143 8483
rect 45143 8449 45152 8483
rect 45100 8440 45152 8449
rect 41972 8372 42024 8424
rect 45468 8508 45520 8560
rect 35072 8347 35124 8356
rect 35072 8313 35081 8347
rect 35081 8313 35115 8347
rect 35115 8313 35124 8347
rect 35072 8304 35124 8313
rect 35808 8347 35860 8356
rect 35808 8313 35817 8347
rect 35817 8313 35851 8347
rect 35851 8313 35860 8347
rect 35808 8304 35860 8313
rect 36452 8304 36504 8356
rect 37004 8304 37056 8356
rect 37096 8304 37148 8356
rect 38752 8347 38804 8356
rect 38752 8313 38761 8347
rect 38761 8313 38795 8347
rect 38795 8313 38804 8347
rect 38752 8304 38804 8313
rect 40132 8304 40184 8356
rect 41604 8304 41656 8356
rect 28172 8236 28224 8288
rect 28540 8236 28592 8288
rect 29184 8279 29236 8288
rect 29184 8245 29193 8279
rect 29193 8245 29227 8279
rect 29227 8245 29236 8279
rect 29184 8236 29236 8245
rect 29276 8236 29328 8288
rect 29920 8279 29972 8288
rect 29920 8245 29929 8279
rect 29929 8245 29963 8279
rect 29963 8245 29972 8279
rect 29920 8236 29972 8245
rect 30288 8279 30340 8288
rect 30288 8245 30297 8279
rect 30297 8245 30331 8279
rect 30331 8245 30340 8279
rect 30288 8236 30340 8245
rect 30380 8236 30432 8288
rect 31392 8279 31444 8288
rect 31392 8245 31401 8279
rect 31401 8245 31435 8279
rect 31435 8245 31444 8279
rect 31392 8236 31444 8245
rect 37648 8279 37700 8288
rect 37648 8245 37657 8279
rect 37657 8245 37691 8279
rect 37691 8245 37700 8279
rect 37648 8236 37700 8245
rect 6665 8134 6717 8186
rect 6729 8134 6781 8186
rect 6793 8134 6845 8186
rect 6857 8134 6909 8186
rect 6921 8134 6973 8186
rect 18095 8134 18147 8186
rect 18159 8134 18211 8186
rect 18223 8134 18275 8186
rect 18287 8134 18339 8186
rect 18351 8134 18403 8186
rect 29525 8134 29577 8186
rect 29589 8134 29641 8186
rect 29653 8134 29705 8186
rect 29717 8134 29769 8186
rect 29781 8134 29833 8186
rect 40955 8134 41007 8186
rect 41019 8134 41071 8186
rect 41083 8134 41135 8186
rect 41147 8134 41199 8186
rect 41211 8134 41263 8186
rect 1124 8032 1176 8084
rect 4068 8075 4120 8084
rect 4068 8041 4077 8075
rect 4077 8041 4111 8075
rect 4111 8041 4120 8075
rect 4068 8032 4120 8041
rect 4804 8032 4856 8084
rect 6552 8032 6604 8084
rect 7380 8032 7432 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 10324 8032 10376 8084
rect 11796 8075 11848 8084
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 12900 8032 12952 8084
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 14740 8032 14792 8084
rect 15844 8032 15896 8084
rect 16672 8032 16724 8084
rect 16948 8032 17000 8084
rect 17684 8032 17736 8084
rect 17960 8032 18012 8084
rect 18420 8032 18472 8084
rect 18788 8075 18840 8084
rect 18788 8041 18797 8075
rect 18797 8041 18831 8075
rect 18831 8041 18840 8075
rect 18788 8032 18840 8041
rect 19524 8032 19576 8084
rect 19984 8032 20036 8084
rect 1860 7896 1912 7948
rect 2136 7803 2188 7812
rect 2136 7769 2145 7803
rect 2145 7769 2179 7803
rect 2179 7769 2188 7803
rect 2136 7760 2188 7769
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 16396 7964 16448 8016
rect 20536 8032 20588 8084
rect 20904 8032 20956 8084
rect 21272 8075 21324 8084
rect 21272 8041 21281 8075
rect 21281 8041 21315 8075
rect 21315 8041 21324 8075
rect 21272 8032 21324 8041
rect 21364 8032 21416 8084
rect 22376 8032 22428 8084
rect 4344 7803 4396 7812
rect 4344 7769 4353 7803
rect 4353 7769 4387 7803
rect 4387 7769 4396 7803
rect 4344 7760 4396 7769
rect 6920 7803 6972 7812
rect 6920 7769 6929 7803
rect 6929 7769 6963 7803
rect 6963 7769 6972 7803
rect 6920 7760 6972 7769
rect 10048 7760 10100 7812
rect 18144 7896 18196 7948
rect 13728 7828 13780 7880
rect 14648 7803 14700 7812
rect 14648 7769 14657 7803
rect 14657 7769 14691 7803
rect 14691 7769 14700 7803
rect 14648 7760 14700 7769
rect 14832 7760 14884 7812
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 17960 7871 18012 7880
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 18420 7828 18472 7880
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 18972 7828 19024 7880
rect 19708 7896 19760 7948
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 20444 7896 20496 7948
rect 20076 7871 20128 7880
rect 20076 7837 20085 7871
rect 20085 7837 20119 7871
rect 20119 7837 20128 7871
rect 20076 7828 20128 7837
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 23480 8032 23532 8084
rect 24216 8032 24268 8084
rect 25136 8032 25188 8084
rect 25412 8075 25464 8084
rect 25412 8041 25421 8075
rect 25421 8041 25455 8075
rect 25455 8041 25464 8075
rect 25412 8032 25464 8041
rect 25504 8032 25556 8084
rect 25872 8032 25924 8084
rect 20720 7828 20772 7880
rect 22468 7896 22520 7948
rect 21180 7871 21232 7880
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 21824 7828 21876 7880
rect 22008 7871 22060 7880
rect 22008 7837 22017 7871
rect 22017 7837 22051 7871
rect 22051 7837 22060 7871
rect 22008 7828 22060 7837
rect 22744 7896 22796 7948
rect 22652 7828 22704 7880
rect 22836 7871 22888 7880
rect 22836 7837 22845 7871
rect 22845 7837 22879 7871
rect 22879 7837 22888 7871
rect 22836 7828 22888 7837
rect 23296 7828 23348 7880
rect 23572 7828 23624 7880
rect 25044 7964 25096 8016
rect 15108 7692 15160 7744
rect 16212 7692 16264 7744
rect 19340 7735 19392 7744
rect 19340 7701 19349 7735
rect 19349 7701 19383 7735
rect 19383 7701 19392 7735
rect 19340 7692 19392 7701
rect 19984 7692 20036 7744
rect 20628 7692 20680 7744
rect 21548 7735 21600 7744
rect 21548 7701 21557 7735
rect 21557 7701 21591 7735
rect 21591 7701 21600 7735
rect 21548 7692 21600 7701
rect 22744 7760 22796 7812
rect 24860 7828 24912 7880
rect 25228 7828 25280 7880
rect 25780 7828 25832 7880
rect 27344 8032 27396 8084
rect 27712 8075 27764 8084
rect 27712 8041 27721 8075
rect 27721 8041 27755 8075
rect 27755 8041 27764 8075
rect 27712 8032 27764 8041
rect 28080 8075 28132 8084
rect 28080 8041 28089 8075
rect 28089 8041 28123 8075
rect 28123 8041 28132 8075
rect 28080 8032 28132 8041
rect 28816 8032 28868 8084
rect 29184 8032 29236 8084
rect 29368 8032 29420 8084
rect 29920 8032 29972 8084
rect 40500 8032 40552 8084
rect 42800 8032 42852 8084
rect 43720 8032 43772 8084
rect 46572 8032 46624 8084
rect 26516 8007 26568 8016
rect 26516 7973 26525 8007
rect 26525 7973 26559 8007
rect 26559 7973 26568 8007
rect 26516 7964 26568 7973
rect 27068 8007 27120 8016
rect 27068 7973 27077 8007
rect 27077 7973 27111 8007
rect 27111 7973 27120 8007
rect 27068 7964 27120 7973
rect 44180 8007 44232 8016
rect 44180 7973 44189 8007
rect 44189 7973 44223 8007
rect 44223 7973 44232 8007
rect 44180 7964 44232 7973
rect 26148 7871 26200 7880
rect 26148 7837 26157 7871
rect 26157 7837 26191 7871
rect 26191 7837 26200 7871
rect 26148 7828 26200 7837
rect 26608 7828 26660 7880
rect 26792 7828 26844 7880
rect 27160 7828 27212 7880
rect 27436 7828 27488 7880
rect 27528 7871 27580 7880
rect 27528 7837 27537 7871
rect 27537 7837 27571 7871
rect 27571 7837 27580 7871
rect 27528 7828 27580 7837
rect 28172 7828 28224 7880
rect 28540 7828 28592 7880
rect 29276 7828 29328 7880
rect 30288 7828 30340 7880
rect 40040 7828 40092 7880
rect 22284 7692 22336 7744
rect 22928 7735 22980 7744
rect 22928 7701 22937 7735
rect 22937 7701 22971 7735
rect 22971 7701 22980 7735
rect 22928 7692 22980 7701
rect 23204 7735 23256 7744
rect 23204 7701 23213 7735
rect 23213 7701 23247 7735
rect 23247 7701 23256 7735
rect 23204 7692 23256 7701
rect 37096 7760 37148 7812
rect 43260 7803 43312 7812
rect 43260 7769 43269 7803
rect 43269 7769 43303 7803
rect 43303 7769 43312 7803
rect 43260 7760 43312 7769
rect 43996 7803 44048 7812
rect 43996 7769 44005 7803
rect 44005 7769 44039 7803
rect 44039 7769 44048 7803
rect 43996 7760 44048 7769
rect 45100 7803 45152 7812
rect 45100 7769 45109 7803
rect 45109 7769 45143 7803
rect 45143 7769 45152 7803
rect 45100 7760 45152 7769
rect 45836 7760 45888 7812
rect 24584 7692 24636 7744
rect 25136 7735 25188 7744
rect 25136 7701 25145 7735
rect 25145 7701 25179 7735
rect 25179 7701 25188 7735
rect 25136 7692 25188 7701
rect 25964 7735 26016 7744
rect 25964 7701 25973 7735
rect 25973 7701 26007 7735
rect 26007 7701 26016 7735
rect 25964 7692 26016 7701
rect 26240 7735 26292 7744
rect 26240 7701 26249 7735
rect 26249 7701 26283 7735
rect 26283 7701 26292 7735
rect 26240 7692 26292 7701
rect 26792 7735 26844 7744
rect 26792 7701 26801 7735
rect 26801 7701 26835 7735
rect 26835 7701 26844 7735
rect 26792 7692 26844 7701
rect 26884 7692 26936 7744
rect 27620 7692 27672 7744
rect 29184 7735 29236 7744
rect 29184 7701 29193 7735
rect 29193 7701 29227 7735
rect 29227 7701 29236 7735
rect 29184 7692 29236 7701
rect 12380 7590 12432 7642
rect 12444 7590 12496 7642
rect 12508 7590 12560 7642
rect 12572 7590 12624 7642
rect 12636 7590 12688 7642
rect 23810 7590 23862 7642
rect 23874 7590 23926 7642
rect 23938 7590 23990 7642
rect 24002 7590 24054 7642
rect 24066 7590 24118 7642
rect 35240 7590 35292 7642
rect 35304 7590 35356 7642
rect 35368 7590 35420 7642
rect 35432 7590 35484 7642
rect 35496 7590 35548 7642
rect 46670 7590 46722 7642
rect 46734 7590 46786 7642
rect 46798 7590 46850 7642
rect 46862 7590 46914 7642
rect 46926 7590 46978 7642
rect 1492 7531 1544 7540
rect 1492 7497 1501 7531
rect 1501 7497 1535 7531
rect 1535 7497 1544 7531
rect 1492 7488 1544 7497
rect 2136 7488 2188 7540
rect 16396 7488 16448 7540
rect 4804 7420 4856 7472
rect 11060 7420 11112 7472
rect 19984 7488 20036 7540
rect 20168 7531 20220 7540
rect 20168 7497 20177 7531
rect 20177 7497 20211 7531
rect 20211 7497 20220 7531
rect 20168 7488 20220 7497
rect 20352 7488 20404 7540
rect 20720 7488 20772 7540
rect 22376 7488 22428 7540
rect 22652 7488 22704 7540
rect 16948 7420 17000 7472
rect 17132 7352 17184 7404
rect 6920 7284 6972 7336
rect 16488 7284 16540 7336
rect 19616 7284 19668 7336
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 20260 7352 20312 7404
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 19708 7216 19760 7268
rect 22560 7352 22612 7404
rect 21180 7284 21232 7336
rect 23296 7488 23348 7540
rect 23388 7488 23440 7540
rect 24768 7488 24820 7540
rect 24860 7488 24912 7540
rect 25044 7488 25096 7540
rect 29000 7488 29052 7540
rect 31392 7488 31444 7540
rect 44548 7488 44600 7540
rect 45284 7488 45336 7540
rect 45652 7531 45704 7540
rect 45652 7497 45661 7531
rect 45661 7497 45695 7531
rect 45695 7497 45704 7531
rect 45652 7488 45704 7497
rect 46388 7531 46440 7540
rect 46388 7497 46397 7531
rect 46397 7497 46431 7531
rect 46431 7497 46440 7531
rect 46388 7488 46440 7497
rect 23480 7352 23532 7404
rect 23664 7352 23716 7404
rect 23848 7395 23900 7404
rect 23848 7361 23857 7395
rect 23857 7361 23891 7395
rect 23891 7361 23900 7395
rect 23848 7352 23900 7361
rect 31116 7420 31168 7472
rect 41604 7352 41656 7404
rect 29092 7284 29144 7336
rect 36452 7284 36504 7336
rect 45560 7395 45612 7404
rect 45560 7361 45569 7395
rect 45569 7361 45603 7395
rect 45603 7361 45612 7395
rect 45560 7352 45612 7361
rect 45652 7352 45704 7404
rect 36912 7216 36964 7268
rect 22744 7148 22796 7200
rect 23388 7191 23440 7200
rect 23388 7157 23397 7191
rect 23397 7157 23431 7191
rect 23431 7157 23440 7191
rect 23388 7148 23440 7157
rect 24032 7191 24084 7200
rect 24032 7157 24041 7191
rect 24041 7157 24075 7191
rect 24075 7157 24084 7191
rect 24032 7148 24084 7157
rect 24676 7148 24728 7200
rect 6665 7046 6717 7098
rect 6729 7046 6781 7098
rect 6793 7046 6845 7098
rect 6857 7046 6909 7098
rect 6921 7046 6973 7098
rect 18095 7046 18147 7098
rect 18159 7046 18211 7098
rect 18223 7046 18275 7098
rect 18287 7046 18339 7098
rect 18351 7046 18403 7098
rect 29525 7046 29577 7098
rect 29589 7046 29641 7098
rect 29653 7046 29705 7098
rect 29717 7046 29769 7098
rect 29781 7046 29833 7098
rect 40955 7046 41007 7098
rect 41019 7046 41071 7098
rect 41083 7046 41135 7098
rect 41147 7046 41199 7098
rect 41211 7046 41263 7098
rect 15752 6944 15804 6996
rect 17040 6944 17092 6996
rect 21180 6944 21232 6996
rect 23480 6944 23532 6996
rect 28908 6944 28960 6996
rect 46020 6944 46072 6996
rect 23388 6876 23440 6928
rect 23848 6876 23900 6928
rect 28448 6876 28500 6928
rect 15292 6808 15344 6860
rect 22928 6808 22980 6860
rect 44916 6808 44968 6860
rect 16120 6740 16172 6792
rect 23204 6740 23256 6792
rect 44364 6740 44416 6792
rect 16488 6672 16540 6724
rect 22652 6672 22704 6724
rect 42800 6672 42852 6724
rect 9680 6604 9732 6656
rect 24032 6604 24084 6656
rect 12380 6502 12432 6554
rect 12444 6502 12496 6554
rect 12508 6502 12560 6554
rect 12572 6502 12624 6554
rect 12636 6502 12688 6554
rect 23810 6502 23862 6554
rect 23874 6502 23926 6554
rect 23938 6502 23990 6554
rect 24002 6502 24054 6554
rect 24066 6502 24118 6554
rect 35240 6502 35292 6554
rect 35304 6502 35356 6554
rect 35368 6502 35420 6554
rect 35432 6502 35484 6554
rect 35496 6502 35548 6554
rect 46670 6502 46722 6554
rect 46734 6502 46786 6554
rect 46798 6502 46850 6554
rect 46862 6502 46914 6554
rect 46926 6502 46978 6554
rect 4344 6400 4396 6452
rect 25136 6400 25188 6452
rect 6460 6332 6512 6384
rect 25964 6332 26016 6384
rect 8300 6264 8352 6316
rect 24584 6264 24636 6316
rect 11060 6196 11112 6248
rect 20720 6196 20772 6248
rect 24768 6128 24820 6180
rect 34520 6128 34572 6180
rect 6665 5958 6717 6010
rect 6729 5958 6781 6010
rect 6793 5958 6845 6010
rect 6857 5958 6909 6010
rect 6921 5958 6973 6010
rect 18095 5958 18147 6010
rect 18159 5958 18211 6010
rect 18223 5958 18275 6010
rect 18287 5958 18339 6010
rect 18351 5958 18403 6010
rect 29525 5958 29577 6010
rect 29589 5958 29641 6010
rect 29653 5958 29705 6010
rect 29717 5958 29769 6010
rect 29781 5958 29833 6010
rect 40955 5958 41007 6010
rect 41019 5958 41071 6010
rect 41083 5958 41135 6010
rect 41147 5958 41199 6010
rect 41211 5958 41263 6010
rect 32128 5584 32180 5636
rect 36636 5584 36688 5636
rect 12380 5414 12432 5466
rect 12444 5414 12496 5466
rect 12508 5414 12560 5466
rect 12572 5414 12624 5466
rect 12636 5414 12688 5466
rect 23810 5414 23862 5466
rect 23874 5414 23926 5466
rect 23938 5414 23990 5466
rect 24002 5414 24054 5466
rect 24066 5414 24118 5466
rect 35240 5414 35292 5466
rect 35304 5414 35356 5466
rect 35368 5414 35420 5466
rect 35432 5414 35484 5466
rect 35496 5414 35548 5466
rect 46670 5414 46722 5466
rect 46734 5414 46786 5466
rect 46798 5414 46850 5466
rect 46862 5414 46914 5466
rect 46926 5414 46978 5466
rect 24676 4972 24728 5024
rect 34612 4972 34664 5024
rect 6665 4870 6717 4922
rect 6729 4870 6781 4922
rect 6793 4870 6845 4922
rect 6857 4870 6909 4922
rect 6921 4870 6973 4922
rect 18095 4870 18147 4922
rect 18159 4870 18211 4922
rect 18223 4870 18275 4922
rect 18287 4870 18339 4922
rect 18351 4870 18403 4922
rect 29525 4870 29577 4922
rect 29589 4870 29641 4922
rect 29653 4870 29705 4922
rect 29717 4870 29769 4922
rect 29781 4870 29833 4922
rect 40955 4870 41007 4922
rect 41019 4870 41071 4922
rect 41083 4870 41135 4922
rect 41147 4870 41199 4922
rect 41211 4870 41263 4922
rect 27712 4768 27764 4820
rect 45100 4768 45152 4820
rect 12380 4326 12432 4378
rect 12444 4326 12496 4378
rect 12508 4326 12560 4378
rect 12572 4326 12624 4378
rect 12636 4326 12688 4378
rect 23810 4326 23862 4378
rect 23874 4326 23926 4378
rect 23938 4326 23990 4378
rect 24002 4326 24054 4378
rect 24066 4326 24118 4378
rect 35240 4326 35292 4378
rect 35304 4326 35356 4378
rect 35368 4326 35420 4378
rect 35432 4326 35484 4378
rect 35496 4326 35548 4378
rect 46670 4326 46722 4378
rect 46734 4326 46786 4378
rect 46798 4326 46850 4378
rect 46862 4326 46914 4378
rect 46926 4326 46978 4378
rect 6665 3782 6717 3834
rect 6729 3782 6781 3834
rect 6793 3782 6845 3834
rect 6857 3782 6909 3834
rect 6921 3782 6973 3834
rect 18095 3782 18147 3834
rect 18159 3782 18211 3834
rect 18223 3782 18275 3834
rect 18287 3782 18339 3834
rect 18351 3782 18403 3834
rect 29525 3782 29577 3834
rect 29589 3782 29641 3834
rect 29653 3782 29705 3834
rect 29717 3782 29769 3834
rect 29781 3782 29833 3834
rect 40955 3782 41007 3834
rect 41019 3782 41071 3834
rect 41083 3782 41135 3834
rect 41147 3782 41199 3834
rect 41211 3782 41263 3834
rect 24216 3612 24268 3664
rect 33692 3612 33744 3664
rect 23664 3544 23716 3596
rect 36084 3544 36136 3596
rect 29920 3476 29972 3528
rect 43996 3476 44048 3528
rect 25688 3408 25740 3460
rect 39948 3408 40000 3460
rect 12380 3238 12432 3290
rect 12444 3238 12496 3290
rect 12508 3238 12560 3290
rect 12572 3238 12624 3290
rect 12636 3238 12688 3290
rect 23810 3238 23862 3290
rect 23874 3238 23926 3290
rect 23938 3238 23990 3290
rect 24002 3238 24054 3290
rect 24066 3238 24118 3290
rect 35240 3238 35292 3290
rect 35304 3238 35356 3290
rect 35368 3238 35420 3290
rect 35432 3238 35484 3290
rect 35496 3238 35548 3290
rect 46670 3238 46722 3290
rect 46734 3238 46786 3290
rect 46798 3238 46850 3290
rect 46862 3238 46914 3290
rect 46926 3238 46978 3290
rect 6665 2694 6717 2746
rect 6729 2694 6781 2746
rect 6793 2694 6845 2746
rect 6857 2694 6909 2746
rect 6921 2694 6973 2746
rect 18095 2694 18147 2746
rect 18159 2694 18211 2746
rect 18223 2694 18275 2746
rect 18287 2694 18339 2746
rect 18351 2694 18403 2746
rect 29525 2694 29577 2746
rect 29589 2694 29641 2746
rect 29653 2694 29705 2746
rect 29717 2694 29769 2746
rect 29781 2694 29833 2746
rect 40955 2694 41007 2746
rect 41019 2694 41071 2746
rect 41083 2694 41135 2746
rect 41147 2694 41199 2746
rect 41211 2694 41263 2746
rect 23664 2635 23716 2644
rect 23664 2601 23673 2635
rect 23673 2601 23707 2635
rect 23707 2601 23716 2635
rect 23664 2592 23716 2601
rect 24216 2635 24268 2644
rect 24216 2601 24225 2635
rect 24225 2601 24259 2635
rect 24259 2601 24268 2635
rect 24216 2592 24268 2601
rect 24768 2635 24820 2644
rect 24768 2601 24777 2635
rect 24777 2601 24811 2635
rect 24811 2601 24820 2635
rect 24768 2592 24820 2601
rect 27620 2592 27672 2644
rect 27712 2635 27764 2644
rect 27712 2601 27721 2635
rect 27721 2601 27755 2635
rect 27755 2601 27764 2635
rect 27712 2592 27764 2601
rect 29920 2635 29972 2644
rect 29920 2601 29929 2635
rect 29929 2601 29963 2635
rect 29963 2601 29972 2635
rect 29920 2592 29972 2601
rect 32128 2635 32180 2644
rect 32128 2601 32137 2635
rect 32137 2601 32171 2635
rect 32171 2601 32180 2635
rect 32128 2592 32180 2601
rect 36452 2592 36504 2644
rect 41604 2592 41656 2644
rect 42800 2592 42852 2644
rect 44364 2592 44416 2644
rect 45560 2592 45612 2644
rect 45652 2635 45704 2644
rect 45652 2601 45661 2635
rect 45661 2601 45695 2635
rect 45695 2601 45704 2635
rect 45652 2592 45704 2601
rect 45744 2635 45796 2644
rect 45744 2601 45753 2635
rect 45753 2601 45787 2635
rect 45787 2601 45796 2635
rect 45744 2592 45796 2601
rect 23480 2524 23532 2576
rect 24768 2456 24820 2508
rect 22376 2388 22428 2440
rect 23664 2388 23716 2440
rect 21088 2363 21140 2372
rect 21088 2329 21097 2363
rect 21097 2329 21131 2363
rect 21131 2329 21140 2363
rect 21088 2320 21140 2329
rect 23204 2363 23256 2372
rect 23204 2329 23213 2363
rect 23213 2329 23247 2363
rect 23247 2329 23256 2363
rect 23204 2320 23256 2329
rect 23572 2320 23624 2372
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 24860 2431 24912 2440
rect 24860 2397 24869 2431
rect 24869 2397 24903 2431
rect 24903 2397 24912 2431
rect 24860 2388 24912 2397
rect 25412 2431 25464 2440
rect 25412 2397 25421 2431
rect 25421 2397 25455 2431
rect 25455 2397 25464 2431
rect 25412 2388 25464 2397
rect 27528 2431 27580 2440
rect 27528 2397 27537 2431
rect 27537 2397 27571 2431
rect 27571 2397 27580 2431
rect 27528 2388 27580 2397
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 31392 2388 31444 2440
rect 34152 2431 34204 2440
rect 34152 2397 34161 2431
rect 34161 2397 34195 2431
rect 34195 2397 34204 2431
rect 34152 2388 34204 2397
rect 40040 2456 40092 2508
rect 40224 2456 40276 2508
rect 36452 2431 36504 2440
rect 36452 2397 36461 2431
rect 36461 2397 36495 2431
rect 36495 2397 36504 2431
rect 36452 2388 36504 2397
rect 38660 2431 38712 2440
rect 38660 2397 38669 2431
rect 38669 2397 38703 2431
rect 38703 2397 38712 2431
rect 38660 2388 38712 2397
rect 43076 2431 43128 2440
rect 43076 2397 43085 2431
rect 43085 2397 43119 2431
rect 43119 2397 43128 2431
rect 43076 2388 43128 2397
rect 45008 2431 45060 2440
rect 45008 2397 45017 2431
rect 45017 2397 45051 2431
rect 45051 2397 45060 2431
rect 45008 2388 45060 2397
rect 21180 2295 21232 2304
rect 21180 2261 21189 2295
rect 21189 2261 21223 2295
rect 21223 2261 21232 2295
rect 21180 2252 21232 2261
rect 24952 2252 25004 2304
rect 33876 2252 33928 2304
rect 40592 2320 40644 2372
rect 44732 2320 44784 2372
rect 45928 2431 45980 2440
rect 45928 2397 45937 2431
rect 45937 2397 45971 2431
rect 45971 2397 45980 2431
rect 45928 2388 45980 2397
rect 12380 2150 12432 2202
rect 12444 2150 12496 2202
rect 12508 2150 12560 2202
rect 12572 2150 12624 2202
rect 12636 2150 12688 2202
rect 23810 2150 23862 2202
rect 23874 2150 23926 2202
rect 23938 2150 23990 2202
rect 24002 2150 24054 2202
rect 24066 2150 24118 2202
rect 35240 2150 35292 2202
rect 35304 2150 35356 2202
rect 35368 2150 35420 2202
rect 35432 2150 35484 2202
rect 35496 2150 35548 2202
rect 46670 2150 46722 2202
rect 46734 2150 46786 2202
rect 46798 2150 46850 2202
rect 46862 2150 46914 2202
rect 46926 2150 46978 2202
rect 21088 2048 21140 2100
rect 21180 2048 21232 2100
rect 22376 2091 22428 2100
rect 22376 2057 22385 2091
rect 22385 2057 22419 2091
rect 22419 2057 22428 2091
rect 22376 2048 22428 2057
rect 23204 2048 23256 2100
rect 23480 2048 23532 2100
rect 24584 2048 24636 2100
rect 25412 2048 25464 2100
rect 27528 2048 27580 2100
rect 29736 2048 29788 2100
rect 31392 2091 31444 2100
rect 31392 2057 31401 2091
rect 31401 2057 31435 2091
rect 31435 2057 31444 2091
rect 31392 2048 31444 2057
rect 34152 2048 34204 2100
rect 36452 2048 36504 2100
rect 38660 2048 38712 2100
rect 43076 2048 43128 2100
rect 43260 2048 43312 2100
rect 45008 2048 45060 2100
rect 45928 2048 45980 2100
rect 20076 1955 20128 1964
rect 20076 1921 20085 1955
rect 20085 1921 20119 1955
rect 20119 1921 20128 1955
rect 20076 1912 20128 1921
rect 20904 1912 20956 1964
rect 22468 1955 22520 1964
rect 22468 1921 22477 1955
rect 22477 1921 22511 1955
rect 22511 1921 22520 1955
rect 22468 1912 22520 1921
rect 22928 1955 22980 1964
rect 22928 1921 22937 1955
rect 22937 1921 22971 1955
rect 22971 1921 22980 1955
rect 22928 1912 22980 1921
rect 19892 1844 19944 1896
rect 23480 1955 23532 1964
rect 23480 1921 23489 1955
rect 23489 1921 23523 1955
rect 23523 1921 23532 1955
rect 23480 1912 23532 1921
rect 23296 1844 23348 1896
rect 24032 1955 24084 1964
rect 24032 1921 24041 1955
rect 24041 1921 24075 1955
rect 24075 1921 24084 1955
rect 24032 1912 24084 1921
rect 24492 1955 24544 1964
rect 24492 1921 24501 1955
rect 24501 1921 24535 1955
rect 24535 1921 24544 1955
rect 24492 1912 24544 1921
rect 24768 1955 24820 1964
rect 24768 1921 24777 1955
rect 24777 1921 24811 1955
rect 24811 1921 24820 1955
rect 24768 1912 24820 1921
rect 24860 1912 24912 1964
rect 26976 1955 27028 1964
rect 26976 1921 26985 1955
rect 26985 1921 27019 1955
rect 27019 1921 27028 1955
rect 26976 1912 27028 1921
rect 29092 1955 29144 1964
rect 29092 1921 29101 1955
rect 29101 1921 29135 1955
rect 29135 1921 29144 1955
rect 29092 1912 29144 1921
rect 31208 1955 31260 1964
rect 31208 1921 31217 1955
rect 31217 1921 31251 1955
rect 31251 1921 31260 1955
rect 31208 1912 31260 1921
rect 33508 1955 33560 1964
rect 33508 1921 33517 1955
rect 33517 1921 33551 1955
rect 33551 1921 33560 1955
rect 33508 1912 33560 1921
rect 35532 1955 35584 1964
rect 35532 1921 35541 1955
rect 35541 1921 35575 1955
rect 35575 1921 35584 1955
rect 35532 1912 35584 1921
rect 37740 1955 37792 1964
rect 37740 1921 37749 1955
rect 37749 1921 37783 1955
rect 37783 1921 37792 1955
rect 37740 1912 37792 1921
rect 42432 1955 42484 1964
rect 42432 1921 42441 1955
rect 42441 1921 42475 1955
rect 42475 1921 42484 1955
rect 42432 1912 42484 1921
rect 44088 1955 44140 1964
rect 44088 1921 44097 1955
rect 44097 1921 44131 1955
rect 44131 1921 44140 1955
rect 44088 1912 44140 1921
rect 44548 1955 44600 1964
rect 44548 1921 44557 1955
rect 44557 1921 44591 1955
rect 44591 1921 44600 1955
rect 44548 1912 44600 1921
rect 45652 1955 45704 1964
rect 45652 1921 45661 1955
rect 45661 1921 45695 1955
rect 45695 1921 45704 1955
rect 45652 1912 45704 1921
rect 23756 1776 23808 1828
rect 25688 1776 25740 1828
rect 44732 1819 44784 1828
rect 44732 1785 44741 1819
rect 44741 1785 44775 1819
rect 44775 1785 44784 1819
rect 44732 1776 44784 1785
rect 24676 1708 24728 1760
rect 27620 1708 27672 1760
rect 36820 1708 36872 1760
rect 6665 1606 6717 1658
rect 6729 1606 6781 1658
rect 6793 1606 6845 1658
rect 6857 1606 6909 1658
rect 6921 1606 6973 1658
rect 18095 1606 18147 1658
rect 18159 1606 18211 1658
rect 18223 1606 18275 1658
rect 18287 1606 18339 1658
rect 18351 1606 18403 1658
rect 29525 1606 29577 1658
rect 29589 1606 29641 1658
rect 29653 1606 29705 1658
rect 29717 1606 29769 1658
rect 29781 1606 29833 1658
rect 40955 1606 41007 1658
rect 41019 1606 41071 1658
rect 41083 1606 41135 1658
rect 41147 1606 41199 1658
rect 41211 1606 41263 1658
rect 20076 1504 20128 1556
rect 22468 1504 22520 1556
rect 23572 1504 23624 1556
rect 24032 1504 24084 1556
rect 24492 1504 24544 1556
rect 26976 1504 27028 1556
rect 29092 1504 29144 1556
rect 31208 1504 31260 1556
rect 33508 1504 33560 1556
rect 35532 1504 35584 1556
rect 37740 1504 37792 1556
rect 42432 1504 42484 1556
rect 44548 1504 44600 1556
rect 45652 1504 45704 1556
rect 15384 1479 15436 1488
rect 15384 1445 15393 1479
rect 15393 1445 15427 1479
rect 15427 1445 15436 1479
rect 15384 1436 15436 1445
rect 1952 1343 2004 1352
rect 1952 1309 1961 1343
rect 1961 1309 1995 1343
rect 1995 1309 2004 1343
rect 1952 1300 2004 1309
rect 4160 1343 4212 1352
rect 4160 1309 4169 1343
rect 4169 1309 4203 1343
rect 4203 1309 4212 1343
rect 4160 1300 4212 1309
rect 6368 1343 6420 1352
rect 6368 1309 6377 1343
rect 6377 1309 6411 1343
rect 6411 1309 6420 1343
rect 6368 1300 6420 1309
rect 8576 1343 8628 1352
rect 8576 1309 8585 1343
rect 8585 1309 8619 1343
rect 8619 1309 8628 1343
rect 8576 1300 8628 1309
rect 10784 1343 10836 1352
rect 10784 1309 10793 1343
rect 10793 1309 10827 1343
rect 10827 1309 10836 1343
rect 10784 1300 10836 1309
rect 12992 1343 13044 1352
rect 12992 1309 13001 1343
rect 13001 1309 13035 1343
rect 13035 1309 13044 1343
rect 12992 1300 13044 1309
rect 15200 1343 15252 1352
rect 15200 1309 15209 1343
rect 15209 1309 15243 1343
rect 15243 1309 15252 1343
rect 15200 1300 15252 1309
rect 17408 1343 17460 1352
rect 17408 1309 17417 1343
rect 17417 1309 17451 1343
rect 17451 1309 17460 1343
rect 17408 1300 17460 1309
rect 19616 1343 19668 1352
rect 19616 1309 19625 1343
rect 19625 1309 19659 1343
rect 19659 1309 19668 1343
rect 19616 1300 19668 1309
rect 2136 1207 2188 1216
rect 2136 1173 2145 1207
rect 2145 1173 2179 1207
rect 2179 1173 2188 1207
rect 2136 1164 2188 1173
rect 20904 1232 20956 1284
rect 6552 1207 6604 1216
rect 6552 1173 6561 1207
rect 6561 1173 6595 1207
rect 6595 1173 6604 1207
rect 6552 1164 6604 1173
rect 8760 1207 8812 1216
rect 8760 1173 8769 1207
rect 8769 1173 8803 1207
rect 8803 1173 8812 1207
rect 8760 1164 8812 1173
rect 10968 1207 11020 1216
rect 10968 1173 10977 1207
rect 10977 1173 11011 1207
rect 11011 1173 11020 1207
rect 10968 1164 11020 1173
rect 15476 1164 15528 1216
rect 21824 1343 21876 1352
rect 21824 1309 21833 1343
rect 21833 1309 21867 1343
rect 21867 1309 21876 1343
rect 21824 1300 21876 1309
rect 23204 1343 23256 1352
rect 23204 1309 23213 1343
rect 23213 1309 23247 1343
rect 23247 1309 23256 1343
rect 23204 1300 23256 1309
rect 21180 1232 21232 1284
rect 24032 1343 24084 1352
rect 24032 1309 24041 1343
rect 24041 1309 24075 1343
rect 24075 1309 24084 1343
rect 24032 1300 24084 1309
rect 26240 1343 26292 1352
rect 26240 1309 26249 1343
rect 26249 1309 26283 1343
rect 26283 1309 26292 1343
rect 26240 1300 26292 1309
rect 28448 1343 28500 1352
rect 28448 1309 28457 1343
rect 28457 1309 28491 1343
rect 28491 1309 28500 1343
rect 28448 1300 28500 1309
rect 30656 1343 30708 1352
rect 30656 1309 30665 1343
rect 30665 1309 30699 1343
rect 30699 1309 30708 1343
rect 30656 1300 30708 1309
rect 32864 1343 32916 1352
rect 32864 1309 32873 1343
rect 32873 1309 32907 1343
rect 32907 1309 32916 1343
rect 32864 1300 32916 1309
rect 35072 1343 35124 1352
rect 35072 1309 35081 1343
rect 35081 1309 35115 1343
rect 35115 1309 35124 1343
rect 35072 1300 35124 1309
rect 37280 1343 37332 1352
rect 37280 1309 37289 1343
rect 37289 1309 37323 1343
rect 37323 1309 37332 1343
rect 37280 1300 37332 1309
rect 39488 1343 39540 1352
rect 39488 1309 39497 1343
rect 39497 1309 39531 1343
rect 39531 1309 39540 1343
rect 39488 1300 39540 1309
rect 41696 1343 41748 1352
rect 41696 1309 41705 1343
rect 41705 1309 41739 1343
rect 41739 1309 41748 1343
rect 41696 1300 41748 1309
rect 43904 1343 43956 1352
rect 43904 1309 43913 1343
rect 43913 1309 43947 1343
rect 43947 1309 43956 1343
rect 43904 1300 43956 1309
rect 46296 1343 46348 1352
rect 46296 1309 46305 1343
rect 46305 1309 46339 1343
rect 46339 1309 46348 1343
rect 46296 1300 46348 1309
rect 23480 1164 23532 1216
rect 44088 1164 44140 1216
rect 12380 1062 12432 1114
rect 12444 1062 12496 1114
rect 12508 1062 12560 1114
rect 12572 1062 12624 1114
rect 12636 1062 12688 1114
rect 23810 1062 23862 1114
rect 23874 1062 23926 1114
rect 23938 1062 23990 1114
rect 24002 1062 24054 1114
rect 24066 1062 24118 1114
rect 35240 1062 35292 1114
rect 35304 1062 35356 1114
rect 35368 1062 35420 1114
rect 35432 1062 35484 1114
rect 35496 1062 35548 1114
rect 46670 1062 46722 1114
rect 46734 1062 46786 1114
rect 46798 1062 46850 1114
rect 46862 1062 46914 1114
rect 46926 1062 46978 1114
rect 2136 960 2188 1012
rect 6552 892 6604 944
rect 8760 960 8812 1012
rect 19892 960 19944 1012
rect 21180 960 21232 1012
rect 23204 960 23256 1012
rect 15384 892 15436 944
rect 15476 892 15528 944
rect 24768 756 24820 808
rect 10968 688 11020 740
rect 23296 688 23348 740
rect 22928 620 22980 672
<< metal2 >>
rect 1122 9840 1178 10000
rect 1490 9840 1546 10000
rect 1858 9840 1914 10000
rect 2226 9840 2282 10000
rect 2594 9840 2650 10000
rect 2962 9840 3018 10000
rect 3330 9840 3386 10000
rect 3698 9840 3754 10000
rect 4066 9840 4122 10000
rect 4434 9840 4490 10000
rect 4802 9840 4858 10000
rect 4908 9846 5120 9874
rect 1136 8090 1164 9840
rect 1124 8084 1176 8090
rect 1124 8026 1176 8032
rect 1504 7546 1532 9840
rect 1872 7954 1900 9840
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8498 1992 8774
rect 2240 8634 2268 9840
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 2332 7857 2360 8434
rect 2608 8430 2636 9840
rect 2976 8634 3004 9840
rect 3344 8634 3372 9840
rect 3712 8634 3740 9840
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2318 7848 2374 7857
rect 2136 7812 2188 7818
rect 2318 7783 2374 7792
rect 2136 7754 2188 7760
rect 2148 7546 2176 7754
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 3252 6905 3280 8434
rect 4080 8090 4108 9840
rect 4448 8634 4476 9840
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4724 8498 4752 8774
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4816 8090 4844 9840
rect 4908 8634 4936 9846
rect 5092 9840 5120 9846
rect 5170 9840 5226 10000
rect 5538 9840 5594 10000
rect 5906 9840 5962 10000
rect 6274 9840 6330 10000
rect 6642 9840 6698 10000
rect 6748 9846 6960 9874
rect 5092 9812 5212 9840
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 5000 8634 5028 9046
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5368 8566 5396 9114
rect 5552 8650 5580 9840
rect 5460 8634 5580 8650
rect 5920 8634 5948 9840
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 5448 8628 5580 8634
rect 5500 8622 5580 8628
rect 5908 8628 5960 8634
rect 5448 8570 5500 8576
rect 5908 8570 5960 8576
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 6196 8498 6224 9590
rect 6288 8634 6316 9840
rect 6656 8786 6684 9840
rect 6564 8758 6684 8786
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 3238 6896 3294 6905
rect 3238 6831 3294 6840
rect 4356 6458 4384 7754
rect 4816 7478 4844 7822
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 6472 6390 6500 8298
rect 6564 8090 6592 8758
rect 6748 8634 6776 9846
rect 6932 9840 6960 9846
rect 7010 9840 7066 10000
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 6932 9812 7052 9840
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 7208 8498 7236 9930
rect 7378 9840 7434 10000
rect 7746 9840 7802 10000
rect 7852 9846 8064 9874
rect 7288 9240 7340 9246
rect 7288 9182 7340 9188
rect 7300 8498 7328 9182
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6665 8188 6973 8197
rect 6665 8186 6671 8188
rect 6727 8186 6751 8188
rect 6807 8186 6831 8188
rect 6887 8186 6911 8188
rect 6967 8186 6973 8188
rect 6727 8134 6729 8186
rect 6909 8134 6911 8186
rect 6665 8132 6671 8134
rect 6727 8132 6751 8134
rect 6807 8132 6831 8134
rect 6887 8132 6911 8134
rect 6967 8132 6973 8134
rect 6665 8123 6973 8132
rect 7392 8090 7420 9840
rect 7760 8634 7788 9840
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7852 8362 7880 9846
rect 8036 9840 8064 9846
rect 8114 9840 8170 10000
rect 8220 9846 8432 9874
rect 8036 9812 8156 9840
rect 8220 8634 8248 9846
rect 8404 9840 8432 9846
rect 8482 9840 8538 10000
rect 8850 9840 8906 10000
rect 9218 9840 9274 10000
rect 9586 9840 9642 10000
rect 9692 9846 9904 9874
rect 8404 9812 8524 9840
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8496 8634 8524 8842
rect 8864 8634 8892 9840
rect 9128 9240 9180 9246
rect 9128 9182 9180 9188
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9140 8498 9168 9182
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 7932 8424 7984 8430
rect 7984 8384 8064 8412
rect 7932 8366 7984 8372
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 8036 8242 8064 8384
rect 8036 8214 8340 8242
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7342 6960 7754
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6665 7100 6973 7109
rect 6665 7098 6671 7100
rect 6727 7098 6751 7100
rect 6807 7098 6831 7100
rect 6887 7098 6911 7100
rect 6967 7098 6973 7100
rect 6727 7046 6729 7098
rect 6909 7046 6911 7098
rect 6665 7044 6671 7046
rect 6727 7044 6751 7046
rect 6807 7044 6831 7046
rect 6887 7044 6911 7046
rect 6967 7044 6973 7046
rect 6665 7035 6973 7044
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 8312 6322 8340 8214
rect 9232 8090 9260 9840
rect 9600 9194 9628 9840
rect 9508 9166 9628 9194
rect 9508 8634 9536 9166
rect 9692 9058 9720 9846
rect 9876 9840 9904 9846
rect 9954 9840 10010 10000
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9876 9812 9996 9840
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 9600 9030 9720 9058
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9600 8566 9628 9030
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9692 6662 9720 8774
rect 10060 8498 10088 9590
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10152 7970 10180 9862
rect 10322 9840 10378 10000
rect 10428 9846 10640 9874
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10244 8498 10272 8978
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10336 8090 10364 9840
rect 10428 8634 10456 9846
rect 10612 9840 10640 9846
rect 10690 9840 10746 10000
rect 11058 9840 11114 10000
rect 11426 9840 11482 10000
rect 11794 9840 11850 10000
rect 12162 9840 12218 10000
rect 12268 9846 12480 9874
rect 10612 9812 10732 9840
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10520 8566 10548 8910
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10612 8498 10640 8774
rect 11072 8650 11100 9840
rect 10980 8634 11100 8650
rect 11440 8634 11468 9840
rect 10968 8628 11100 8634
rect 11020 8622 11100 8628
rect 11428 8628 11480 8634
rect 10968 8570 11020 8576
rect 11428 8570 11480 8576
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 11808 8090 11836 9840
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11900 8498 11928 9658
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11992 8265 12020 9114
rect 12084 8974 12112 9114
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12176 8634 12204 9840
rect 12268 8634 12296 9846
rect 12452 9738 12480 9846
rect 12530 9840 12586 10000
rect 12716 9852 12768 9858
rect 12544 9738 12572 9840
rect 12898 9840 12954 10000
rect 13266 9840 13322 10000
rect 13634 9840 13690 10000
rect 14002 9840 14058 10000
rect 14370 9840 14426 10000
rect 14738 9840 14794 10000
rect 15106 9840 15162 10000
rect 15474 9840 15530 10000
rect 15842 9840 15898 10000
rect 16120 9852 16172 9858
rect 12716 9794 12768 9800
rect 12452 9710 12572 9738
rect 12728 9450 12756 9794
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12380 8732 12688 8741
rect 12380 8730 12386 8732
rect 12442 8730 12466 8732
rect 12522 8730 12546 8732
rect 12602 8730 12626 8732
rect 12682 8730 12688 8732
rect 12442 8678 12444 8730
rect 12624 8678 12626 8730
rect 12380 8676 12386 8678
rect 12442 8676 12466 8678
rect 12522 8676 12546 8678
rect 12602 8676 12626 8678
rect 12682 8676 12688 8678
rect 12380 8667 12688 8676
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12820 8498 12848 9386
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 11978 8256 12034 8265
rect 11978 8191 12034 8200
rect 12912 8090 12940 9840
rect 12990 9072 13046 9081
rect 12990 9007 13046 9016
rect 13004 8498 13032 9007
rect 13280 8634 13308 9840
rect 13648 9432 13676 9840
rect 13464 9404 13676 9432
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8498 13400 8842
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13464 8362 13492 9404
rect 13636 9308 13688 9314
rect 13636 9250 13688 9256
rect 13648 9042 13676 9250
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13726 8936 13782 8945
rect 13544 8900 13596 8906
rect 13726 8871 13782 8880
rect 13544 8842 13596 8848
rect 13556 8498 13584 8842
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 10060 7942 10180 7970
rect 10060 7818 10088 7942
rect 13740 7886 13768 8871
rect 14016 8634 14044 9840
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14384 8090 14412 9840
rect 14646 9208 14702 9217
rect 14646 9143 14702 9152
rect 14660 8498 14688 9143
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14462 8392 14518 8401
rect 14462 8327 14464 8336
rect 14516 8327 14518 8336
rect 14464 8298 14516 8304
rect 14752 8090 14780 9840
rect 15120 8650 15148 9840
rect 14936 8634 15148 8650
rect 15488 8634 15516 9840
rect 14924 8628 15148 8634
rect 14976 8622 15148 8628
rect 15476 8628 15528 8634
rect 14924 8570 14976 8576
rect 15476 8570 15528 8576
rect 14832 8560 14884 8566
rect 14830 8528 14832 8537
rect 14884 8528 14886 8537
rect 14830 8463 14886 8472
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 12380 7644 12688 7653
rect 12380 7642 12386 7644
rect 12442 7642 12466 7644
rect 12522 7642 12546 7644
rect 12602 7642 12626 7644
rect 12682 7642 12688 7644
rect 12442 7590 12444 7642
rect 12624 7590 12626 7642
rect 12380 7588 12386 7590
rect 12442 7588 12466 7590
rect 12522 7588 12546 7590
rect 12602 7588 12626 7590
rect 12682 7588 12688 7590
rect 12380 7579 12688 7588
rect 14660 7585 14688 7754
rect 14646 7576 14702 7585
rect 14646 7511 14702 7520
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 11072 6254 11100 7414
rect 14844 7313 14872 7754
rect 15108 7744 15160 7750
rect 15106 7712 15108 7721
rect 15160 7712 15162 7721
rect 15106 7647 15162 7656
rect 14830 7304 14886 7313
rect 14830 7239 14886 7248
rect 15304 6866 15332 8434
rect 15856 8090 15884 9840
rect 16210 9840 16266 10000
rect 16578 9840 16634 10000
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16120 9794 16172 9800
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7002 15792 7822
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 16132 6798 16160 9794
rect 16224 8634 16252 9840
rect 16592 8650 16620 9840
rect 16868 9625 16896 9930
rect 16946 9840 17002 10000
rect 17314 9840 17370 10000
rect 17682 9840 17738 10000
rect 18050 9840 18106 10000
rect 18418 9840 18474 10000
rect 18786 9840 18842 10000
rect 19154 9840 19210 10000
rect 19522 9840 19578 10000
rect 19890 9840 19946 10000
rect 20258 9840 20314 10000
rect 20626 9840 20682 10000
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 16854 9616 16910 9625
rect 16854 9551 16910 9560
rect 16500 8634 16620 8650
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16488 8628 16620 8634
rect 16540 8622 16620 8628
rect 16488 8570 16540 8576
rect 16210 8256 16266 8265
rect 16210 8191 16266 8200
rect 16224 7750 16252 8191
rect 16960 8090 16988 9840
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17144 9489 17172 9522
rect 17130 9480 17186 9489
rect 17130 9415 17186 9424
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16396 8016 16448 8022
rect 16396 7958 16448 7964
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16408 7546 16436 7958
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16684 7449 16712 8026
rect 16946 7576 17002 7585
rect 16946 7511 17002 7520
rect 16960 7478 16988 7511
rect 16948 7472 17000 7478
rect 16670 7440 16726 7449
rect 16948 7414 17000 7420
rect 16670 7375 16726 7384
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16500 6730 16528 7278
rect 17052 7002 17080 8434
rect 17144 7410 17172 8502
rect 17236 8498 17264 9046
rect 17328 8634 17356 9840
rect 17408 9784 17460 9790
rect 17408 9726 17460 9732
rect 17420 9450 17448 9726
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17696 8634 17724 9840
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17788 9081 17816 9590
rect 17880 9217 17908 9658
rect 17866 9208 17922 9217
rect 17866 9143 17922 9152
rect 17774 9072 17830 9081
rect 17774 9007 17830 9016
rect 18064 8634 18092 9840
rect 18432 8634 18460 9840
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17236 7886 17264 8298
rect 17696 8090 17724 8434
rect 17972 8090 18000 8434
rect 18095 8188 18403 8197
rect 18095 8186 18101 8188
rect 18157 8186 18181 8188
rect 18237 8186 18261 8188
rect 18317 8186 18341 8188
rect 18397 8186 18403 8188
rect 18157 8134 18159 8186
rect 18339 8134 18341 8186
rect 18095 8132 18101 8134
rect 18157 8132 18181 8134
rect 18237 8132 18261 8134
rect 18317 8132 18341 8134
rect 18397 8132 18403 8134
rect 18095 8123 18403 8132
rect 18432 8090 18460 8434
rect 18510 8120 18566 8129
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18420 8084 18472 8090
rect 18510 8055 18566 8064
rect 18420 8026 18472 8032
rect 17958 7984 18014 7993
rect 17958 7919 18014 7928
rect 18144 7948 18196 7954
rect 17972 7886 18000 7919
rect 18144 7890 18196 7896
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18156 7585 18184 7890
rect 18524 7886 18552 8055
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18432 7732 18460 7822
rect 18616 7732 18644 9454
rect 18800 8634 18828 9840
rect 18970 9752 19026 9761
rect 18970 9687 19026 9696
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18800 8090 18828 8434
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18984 7886 19012 9687
rect 19062 9616 19118 9625
rect 19062 9551 19118 9560
rect 19076 8378 19104 9551
rect 19168 9058 19196 9840
rect 19168 9030 19288 9058
rect 19260 8566 19288 9030
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19536 8430 19564 9840
rect 19798 9344 19854 9353
rect 19798 9279 19854 9288
rect 19706 8664 19762 8673
rect 19706 8599 19762 8608
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19524 8424 19576 8430
rect 19076 8350 19288 8378
rect 19524 8366 19576 8372
rect 19260 8242 19288 8350
rect 19338 8256 19394 8265
rect 19260 8214 19338 8242
rect 19338 8191 19394 8200
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19536 7886 19564 8026
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 18432 7704 18644 7732
rect 19340 7744 19392 7750
rect 19338 7712 19340 7721
rect 19392 7712 19394 7721
rect 19338 7647 19394 7656
rect 18142 7576 18198 7585
rect 18142 7511 18198 7520
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 19628 7342 19656 8434
rect 19720 8362 19748 8599
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19720 7274 19748 7890
rect 19812 7410 19840 9279
rect 19904 8634 19932 9840
rect 19984 9648 20036 9654
rect 19982 9616 19984 9625
rect 20036 9616 20038 9625
rect 19982 9551 20038 9560
rect 20074 9208 20130 9217
rect 20074 9143 20130 9152
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19996 8090 20024 8434
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 20088 7886 20116 9143
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19996 7546 20024 7686
rect 20180 7546 20208 8434
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20272 7410 20300 9840
rect 20352 9104 20404 9110
rect 20352 9046 20404 9052
rect 20364 8634 20392 9046
rect 20640 8922 20668 9840
rect 20456 8894 20668 8922
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20456 7954 20484 8894
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20548 8090 20576 8570
rect 20732 8378 20760 9862
rect 20916 9625 20944 9862
rect 20994 9840 21050 10000
rect 21100 9846 21312 9874
rect 20902 9616 20958 9625
rect 20902 9551 20958 9560
rect 21008 8650 21036 9840
rect 20640 8350 20760 8378
rect 20824 8622 21036 8650
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 7546 20392 7822
rect 20640 7750 20668 8350
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20732 7886 20760 8230
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19996 7177 20024 7346
rect 19982 7168 20038 7177
rect 18095 7100 18403 7109
rect 19982 7103 20038 7112
rect 18095 7098 18101 7100
rect 18157 7098 18181 7100
rect 18237 7098 18261 7100
rect 18317 7098 18341 7100
rect 18397 7098 18403 7100
rect 18157 7046 18159 7098
rect 18339 7046 18341 7098
rect 18095 7044 18101 7046
rect 18157 7044 18181 7046
rect 18237 7044 18261 7046
rect 18317 7044 18341 7046
rect 18397 7044 18403 7046
rect 18095 7035 18403 7044
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 12380 6556 12688 6565
rect 12380 6554 12386 6556
rect 12442 6554 12466 6556
rect 12522 6554 12546 6556
rect 12602 6554 12626 6556
rect 12682 6554 12688 6556
rect 12442 6502 12444 6554
rect 12624 6502 12626 6554
rect 12380 6500 12386 6502
rect 12442 6500 12466 6502
rect 12522 6500 12546 6502
rect 12602 6500 12626 6502
rect 12682 6500 12688 6502
rect 12380 6491 12688 6500
rect 20732 6254 20760 7482
rect 20824 7410 20852 8622
rect 21100 8498 21128 9846
rect 21284 9738 21312 9846
rect 21362 9840 21418 10000
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21376 9738 21404 9840
rect 21284 9710 21404 9738
rect 21178 9480 21234 9489
rect 21234 9438 21312 9466
rect 21178 9415 21234 9424
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 20902 8392 20958 8401
rect 20902 8327 20958 8336
rect 20916 8090 20944 8327
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 21192 7886 21220 8230
rect 21284 8090 21312 9438
rect 21364 9240 21416 9246
rect 21364 9182 21416 9188
rect 21456 9240 21508 9246
rect 21456 9182 21508 9188
rect 21376 8809 21404 9182
rect 21362 8800 21418 8809
rect 21362 8735 21418 8744
rect 21468 8634 21496 9182
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21560 8401 21588 9930
rect 21730 9840 21786 10000
rect 22098 9840 22154 10000
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22192 9852 22244 9858
rect 21638 9752 21694 9761
rect 21638 9687 21694 9696
rect 21652 9178 21680 9687
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21638 9072 21694 9081
rect 21638 9007 21640 9016
rect 21692 9007 21694 9016
rect 21640 8978 21692 8984
rect 21744 8566 21772 9840
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21836 9353 21864 9454
rect 21822 9344 21878 9353
rect 21822 9279 21878 9288
rect 22020 8906 22048 9454
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21824 8492 21876 8498
rect 22112 8480 22140 9840
rect 22192 9794 22244 9800
rect 22204 9654 22232 9794
rect 22192 9648 22244 9654
rect 22296 9625 22324 9862
rect 22466 9840 22522 10000
rect 22572 9846 22784 9874
rect 22192 9590 22244 9596
rect 22282 9616 22338 9625
rect 22480 9568 22508 9840
rect 22282 9551 22338 9560
rect 22388 9540 22508 9568
rect 22388 9432 22416 9540
rect 22296 9404 22416 9432
rect 22192 9240 22244 9246
rect 22192 9182 22244 9188
rect 21876 8452 22140 8480
rect 21824 8434 21876 8440
rect 21546 8392 21602 8401
rect 22204 8378 22232 9182
rect 22296 8634 22324 9404
rect 22376 9308 22428 9314
rect 22376 9250 22428 9256
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 22204 8362 22324 8378
rect 22204 8356 22336 8362
rect 22204 8350 22284 8356
rect 21546 8327 21602 8336
rect 22284 8298 22336 8304
rect 21456 8288 21508 8294
rect 21362 8256 21418 8265
rect 21456 8230 21508 8236
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 22008 8288 22060 8294
rect 22388 8242 22416 9250
rect 22468 9104 22520 9110
rect 22466 9072 22468 9081
rect 22520 9072 22522 9081
rect 22466 9007 22522 9016
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22008 8230 22060 8236
rect 21362 8191 21418 8200
rect 21376 8090 21404 8191
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21468 7886 21496 8230
rect 21836 7886 21864 8230
rect 22020 7886 22048 8230
rect 22296 8214 22416 8242
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 22296 7750 22324 8214
rect 22376 8084 22428 8090
rect 22376 8026 22428 8032
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 21560 7585 21588 7686
rect 21546 7576 21602 7585
rect 22388 7546 22416 8026
rect 22480 7954 22508 8842
rect 22572 8634 22600 9846
rect 22756 9840 22784 9846
rect 22834 9840 22890 10000
rect 22940 9846 23152 9874
rect 22756 9812 22876 9840
rect 22650 9752 22706 9761
rect 22650 9687 22652 9696
rect 22704 9687 22706 9696
rect 22652 9658 22704 9664
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22756 8809 22784 8978
rect 22742 8800 22798 8809
rect 22742 8735 22798 8744
rect 22650 8664 22706 8673
rect 22560 8628 22612 8634
rect 22650 8599 22652 8608
rect 22560 8570 22612 8576
rect 22704 8599 22706 8608
rect 22652 8570 22704 8576
rect 22560 8492 22612 8498
rect 22940 8480 22968 9846
rect 23124 9840 23152 9846
rect 23202 9840 23258 10000
rect 23308 9846 23520 9874
rect 23124 9812 23244 9840
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 23032 8634 23060 8774
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 23124 8498 23152 8910
rect 23204 8560 23256 8566
rect 23308 8548 23336 9846
rect 23492 9840 23520 9846
rect 23570 9840 23626 10000
rect 23676 9846 23888 9874
rect 23492 9812 23612 9840
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23256 8520 23336 8548
rect 23204 8502 23256 8508
rect 22612 8452 22968 8480
rect 23112 8492 23164 8498
rect 22560 8434 22612 8440
rect 23112 8434 23164 8440
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22744 8288 22796 8294
rect 22744 8230 22796 8236
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 21546 7511 21602 7520
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22572 7410 22600 8230
rect 22664 7886 22692 8230
rect 22756 7954 22784 8230
rect 23492 8090 23520 9522
rect 23584 8378 23612 9522
rect 23676 8548 23704 9846
rect 23860 9840 23888 9846
rect 23938 9840 23994 10000
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 23860 9812 23980 9840
rect 24044 9353 24072 9930
rect 24306 9840 24362 10000
rect 24400 9852 24452 9858
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24030 9344 24086 9353
rect 24030 9279 24086 9288
rect 24136 8838 24164 9590
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 23810 8732 24118 8741
rect 23810 8730 23816 8732
rect 23872 8730 23896 8732
rect 23952 8730 23976 8732
rect 24032 8730 24056 8732
rect 24112 8730 24118 8732
rect 23872 8678 23874 8730
rect 24054 8678 24056 8730
rect 23810 8676 23816 8678
rect 23872 8676 23896 8678
rect 23952 8676 23976 8678
rect 24032 8676 24056 8678
rect 24112 8676 24118 8678
rect 23810 8667 24118 8676
rect 23756 8560 23808 8566
rect 23676 8520 23756 8548
rect 23756 8502 23808 8508
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23756 8424 23808 8430
rect 23754 8392 23756 8401
rect 23808 8392 23810 8401
rect 23584 8350 23704 8378
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 23584 7886 23612 8230
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 22744 7812 22796 7818
rect 22744 7754 22796 7760
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 21192 7002 21220 7278
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 22664 6730 22692 7482
rect 22756 7206 22784 7754
rect 22848 7721 22876 7822
rect 22928 7744 22980 7750
rect 22834 7712 22890 7721
rect 22928 7686 22980 7692
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 22834 7647 22890 7656
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22940 6866 22968 7686
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 23216 6798 23244 7686
rect 23308 7546 23336 7822
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23400 7449 23428 7482
rect 23386 7440 23442 7449
rect 23676 7410 23704 8350
rect 23754 8327 23810 8336
rect 23860 8265 23888 8434
rect 23846 8256 23902 8265
rect 23846 8191 23902 8200
rect 24228 8090 24256 9658
rect 24320 8566 24348 9840
rect 24674 9840 24730 10000
rect 24780 9846 24992 9874
rect 24780 9840 24808 9846
rect 24688 9812 24808 9840
rect 24400 9794 24452 9800
rect 24412 9586 24440 9794
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24688 9217 24716 9522
rect 24768 9512 24820 9518
rect 24766 9480 24768 9489
rect 24820 9480 24822 9489
rect 24766 9415 24822 9424
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24674 9208 24730 9217
rect 24674 9143 24730 9152
rect 24676 9036 24728 9042
rect 24676 8978 24728 8984
rect 24308 8560 24360 8566
rect 24308 8502 24360 8508
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 24412 8401 24440 8434
rect 24398 8392 24454 8401
rect 24398 8327 24454 8336
rect 24216 8084 24268 8090
rect 24216 8026 24268 8032
rect 24584 7744 24636 7750
rect 24584 7686 24636 7692
rect 23810 7644 24118 7653
rect 23810 7642 23816 7644
rect 23872 7642 23896 7644
rect 23952 7642 23976 7644
rect 24032 7642 24056 7644
rect 24112 7642 24118 7644
rect 23872 7590 23874 7642
rect 24054 7590 24056 7642
rect 23810 7588 23816 7590
rect 23872 7588 23896 7590
rect 23952 7588 23976 7590
rect 24032 7588 24056 7590
rect 24112 7588 24118 7590
rect 23810 7579 24118 7588
rect 23386 7375 23442 7384
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23400 6934 23428 7142
rect 23492 7002 23520 7346
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 23860 6934 23888 7346
rect 24032 7200 24084 7206
rect 24032 7142 24084 7148
rect 23388 6928 23440 6934
rect 23388 6870 23440 6876
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 22652 6724 22704 6730
rect 22652 6666 22704 6672
rect 24044 6662 24072 7142
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 23810 6556 24118 6565
rect 23810 6554 23816 6556
rect 23872 6554 23896 6556
rect 23952 6554 23976 6556
rect 24032 6554 24056 6556
rect 24112 6554 24118 6556
rect 23872 6502 23874 6554
rect 24054 6502 24056 6554
rect 23810 6500 23816 6502
rect 23872 6500 23896 6502
rect 23952 6500 23976 6502
rect 24032 6500 24056 6502
rect 24112 6500 24118 6502
rect 23810 6491 24118 6500
rect 24596 6322 24624 7686
rect 24688 7206 24716 8978
rect 24872 8906 24900 9318
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24964 8498 24992 9846
rect 25042 9840 25098 10000
rect 25148 9846 25360 9874
rect 25148 9840 25176 9846
rect 25056 9812 25176 9840
rect 25332 8498 25360 9846
rect 25410 9840 25466 10000
rect 25516 9846 25728 9874
rect 25516 9840 25544 9846
rect 25424 9812 25544 9840
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25410 8528 25466 8537
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 25320 8492 25372 8498
rect 25410 8463 25466 8472
rect 25320 8434 25372 8440
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 24780 7546 24808 8230
rect 25148 8090 25176 8230
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25044 8016 25096 8022
rect 25044 7958 25096 7964
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24872 7546 24900 7822
rect 25056 7546 25084 7958
rect 25240 7886 25268 8230
rect 25424 8090 25452 8463
rect 25516 8090 25544 9046
rect 25700 8498 25728 9846
rect 25778 9840 25834 10000
rect 25884 9846 26096 9874
rect 25884 9840 25912 9846
rect 25792 9812 25912 9840
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 25504 8084 25556 8090
rect 25504 8026 25556 8032
rect 25792 7886 25820 8570
rect 26068 8498 26096 9846
rect 26146 9840 26202 10000
rect 26252 9846 26464 9874
rect 26252 9840 26280 9846
rect 26160 9812 26280 9840
rect 26436 8498 26464 9846
rect 26514 9840 26570 10000
rect 26620 9846 26832 9874
rect 26620 9840 26648 9846
rect 26528 9812 26648 9840
rect 26516 9444 26568 9450
rect 26516 9386 26568 9392
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26148 8356 26200 8362
rect 26148 8298 26200 8304
rect 25872 8288 25924 8294
rect 25872 8230 25924 8236
rect 25884 8090 25912 8230
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 26160 7886 26188 8298
rect 26528 8022 26556 9386
rect 26804 8498 26832 9846
rect 26882 9840 26938 10000
rect 26988 9846 27200 9874
rect 26988 9840 27016 9846
rect 26896 9812 27016 9840
rect 27068 9784 27120 9790
rect 27068 9726 27120 9732
rect 26884 9240 26936 9246
rect 26884 9182 26936 9188
rect 26792 8492 26844 8498
rect 26792 8434 26844 8440
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26516 8016 26568 8022
rect 26516 7958 26568 7964
rect 26620 7886 26648 8230
rect 26804 7886 26832 8230
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26896 7750 26924 9182
rect 27080 8022 27108 9726
rect 27172 8498 27200 9846
rect 27250 9840 27306 10000
rect 27356 9846 27568 9874
rect 27356 9840 27384 9846
rect 27264 9812 27384 9840
rect 27344 8560 27396 8566
rect 27344 8502 27396 8508
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27160 8288 27212 8294
rect 27160 8230 27212 8236
rect 27068 8016 27120 8022
rect 27068 7958 27120 7964
rect 27172 7886 27200 8230
rect 27356 8090 27384 8502
rect 27540 8498 27568 9846
rect 27618 9840 27674 10000
rect 27724 9846 27936 9874
rect 27724 9840 27752 9846
rect 27632 9812 27752 9840
rect 27710 9616 27766 9625
rect 27710 9551 27766 9560
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 27448 7886 27476 8298
rect 27528 8288 27580 8294
rect 27528 8230 27580 8236
rect 27540 7886 27568 8230
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27632 7750 27660 8774
rect 27724 8090 27752 9551
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27816 8838 27844 9318
rect 27804 8832 27856 8838
rect 27804 8774 27856 8780
rect 27908 8498 27936 9846
rect 27986 9840 28042 10000
rect 28092 9846 28304 9874
rect 28092 9840 28120 9846
rect 28000 9812 28120 9840
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 27712 8084 27764 8090
rect 27712 8026 27764 8032
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 26240 7744 26292 7750
rect 26792 7744 26844 7750
rect 26240 7686 26292 7692
rect 26790 7712 26792 7721
rect 26884 7744 26936 7750
rect 26844 7712 26846 7721
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 25148 6458 25176 7686
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25976 6390 26004 7686
rect 26252 6905 26280 7686
rect 26884 7686 26936 7692
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 26790 7647 26846 7656
rect 28000 7177 28028 9114
rect 28078 8936 28134 8945
rect 28078 8871 28134 8880
rect 28092 8090 28120 8871
rect 28184 8401 28212 9522
rect 28276 8498 28304 9846
rect 28354 9840 28410 10000
rect 28460 9846 28672 9874
rect 28460 9840 28488 9846
rect 28368 9812 28488 9840
rect 28354 9752 28410 9761
rect 28354 9687 28410 9696
rect 28368 9314 28396 9687
rect 28356 9308 28408 9314
rect 28356 9250 28408 9256
rect 28448 9240 28500 9246
rect 28448 9182 28500 9188
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28170 8392 28226 8401
rect 28170 8327 28226 8336
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 28262 8256 28318 8265
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 28184 7886 28212 8230
rect 28368 8242 28396 8910
rect 28318 8214 28396 8242
rect 28262 8191 28318 8200
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 27986 7168 28042 7177
rect 27986 7103 28042 7112
rect 28460 6934 28488 9182
rect 28644 8498 28672 9846
rect 28722 9840 28778 10000
rect 28816 9920 28868 9926
rect 28816 9862 28868 9868
rect 28908 9920 28960 9926
rect 28908 9862 28960 9868
rect 28736 8498 28764 9840
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 28540 8288 28592 8294
rect 28540 8230 28592 8236
rect 28552 7886 28580 8230
rect 28828 8090 28856 9862
rect 28816 8084 28868 8090
rect 28816 8026 28868 8032
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28920 7002 28948 9862
rect 29090 9840 29146 10000
rect 29196 9846 29408 9874
rect 29196 9840 29224 9846
rect 29104 9812 29224 9840
rect 29276 9716 29328 9722
rect 29276 9658 29328 9664
rect 29092 9104 29144 9110
rect 29092 9046 29144 9052
rect 29000 8356 29052 8362
rect 29000 8298 29052 8304
rect 29012 7546 29040 8298
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 29104 7342 29132 9046
rect 29288 8378 29316 9658
rect 29380 8498 29408 9846
rect 29458 9840 29514 10000
rect 29564 9846 29776 9874
rect 29564 9840 29592 9846
rect 29472 9812 29592 9840
rect 29748 8498 29776 9846
rect 29826 9840 29882 10000
rect 29932 9846 30144 9874
rect 29932 9840 29960 9846
rect 29840 9812 29960 9840
rect 30116 8498 30144 9846
rect 30194 9840 30250 10000
rect 30562 9840 30618 10000
rect 30930 9840 30986 10000
rect 31036 9846 31248 9874
rect 31036 9840 31064 9846
rect 30208 8498 30236 9840
rect 30576 8616 30604 9840
rect 30944 9812 31064 9840
rect 30748 8628 30800 8634
rect 30576 8588 30748 8616
rect 30748 8570 30800 8576
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 30380 8560 30432 8566
rect 30380 8502 30432 8508
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 29288 8350 29408 8378
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29276 8288 29328 8294
rect 29276 8230 29328 8236
rect 29196 8090 29224 8230
rect 29184 8084 29236 8090
rect 29184 8026 29236 8032
rect 29288 7886 29316 8230
rect 29380 8090 29408 8350
rect 30392 8294 30420 8502
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 30288 8288 30340 8294
rect 30288 8230 30340 8236
rect 30380 8288 30432 8294
rect 30380 8230 30432 8236
rect 29525 8188 29833 8197
rect 29525 8186 29531 8188
rect 29587 8186 29611 8188
rect 29667 8186 29691 8188
rect 29747 8186 29771 8188
rect 29827 8186 29833 8188
rect 29587 8134 29589 8186
rect 29769 8134 29771 8186
rect 29525 8132 29531 8134
rect 29587 8132 29611 8134
rect 29667 8132 29691 8134
rect 29747 8132 29771 8134
rect 29827 8132 29833 8134
rect 29525 8123 29833 8132
rect 29932 8090 29960 8230
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 30300 7886 30328 8230
rect 29276 7880 29328 7886
rect 29276 7822 29328 7828
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 29184 7744 29236 7750
rect 29184 7686 29236 7692
rect 29092 7336 29144 7342
rect 29196 7313 29224 7686
rect 31128 7478 31156 8570
rect 31220 8498 31248 9846
rect 31298 9840 31354 10000
rect 31404 9846 31616 9874
rect 31404 9840 31432 9846
rect 31312 9812 31432 9840
rect 31588 8498 31616 9846
rect 31666 9840 31722 10000
rect 32034 9840 32090 10000
rect 32140 9846 32352 9874
rect 32140 9840 32168 9846
rect 31680 8498 31708 9840
rect 32048 9812 32168 9840
rect 32128 9104 32180 9110
rect 32128 9046 32180 9052
rect 32140 8634 32168 9046
rect 32128 8628 32180 8634
rect 32128 8570 32180 8576
rect 32324 8498 32352 9846
rect 32402 9840 32458 10000
rect 32508 9846 32720 9874
rect 32508 9840 32536 9846
rect 32416 9812 32536 9840
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 32600 8634 32628 9318
rect 32588 8628 32640 8634
rect 32588 8570 32640 8576
rect 32692 8498 32720 9846
rect 32770 9840 32826 10000
rect 32876 9846 33088 9874
rect 32876 9840 32904 9846
rect 32784 9812 32904 9840
rect 33060 8498 33088 9846
rect 33138 9840 33194 10000
rect 33244 9846 33456 9874
rect 33244 9840 33272 9846
rect 33152 9812 33272 9840
rect 33232 9580 33284 9586
rect 33232 9522 33284 9528
rect 33244 8634 33272 9522
rect 33232 8628 33284 8634
rect 33232 8570 33284 8576
rect 33428 8498 33456 9846
rect 33506 9840 33562 10000
rect 33612 9846 33824 9874
rect 33612 9840 33640 9846
rect 33520 9812 33640 9840
rect 33600 9512 33652 9518
rect 33600 9454 33652 9460
rect 33612 8634 33640 9454
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33796 8498 33824 9846
rect 33874 9840 33930 10000
rect 33980 9846 34192 9874
rect 33980 9840 34008 9846
rect 33888 9812 34008 9840
rect 33876 9376 33928 9382
rect 33876 9318 33928 9324
rect 31208 8492 31260 8498
rect 31208 8434 31260 8440
rect 31576 8492 31628 8498
rect 31576 8434 31628 8440
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 33048 8492 33100 8498
rect 33048 8434 33100 8440
rect 33416 8492 33468 8498
rect 33416 8434 33468 8440
rect 33784 8492 33836 8498
rect 33784 8434 33836 8440
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 31392 8288 31444 8294
rect 31392 8230 31444 8236
rect 31404 7546 31432 8230
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31116 7472 31168 7478
rect 31116 7414 31168 7420
rect 29092 7278 29144 7284
rect 29182 7304 29238 7313
rect 29182 7239 29238 7248
rect 29525 7100 29833 7109
rect 29525 7098 29531 7100
rect 29587 7098 29611 7100
rect 29667 7098 29691 7100
rect 29747 7098 29771 7100
rect 29827 7098 29833 7100
rect 29587 7046 29589 7098
rect 29769 7046 29771 7098
rect 29525 7044 29531 7046
rect 29587 7044 29611 7046
rect 29667 7044 29691 7046
rect 29747 7044 29771 7046
rect 29827 7044 29833 7046
rect 29525 7035 29833 7044
rect 28908 6996 28960 7002
rect 28908 6938 28960 6944
rect 28448 6928 28500 6934
rect 26238 6896 26294 6905
rect 28448 6870 28500 6876
rect 26238 6831 26294 6840
rect 25964 6384 26016 6390
rect 25964 6326 26016 6332
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 6665 6012 6973 6021
rect 6665 6010 6671 6012
rect 6727 6010 6751 6012
rect 6807 6010 6831 6012
rect 6887 6010 6911 6012
rect 6967 6010 6973 6012
rect 6727 5958 6729 6010
rect 6909 5958 6911 6010
rect 6665 5956 6671 5958
rect 6727 5956 6751 5958
rect 6807 5956 6831 5958
rect 6887 5956 6911 5958
rect 6967 5956 6973 5958
rect 6665 5947 6973 5956
rect 18095 6012 18403 6021
rect 18095 6010 18101 6012
rect 18157 6010 18181 6012
rect 18237 6010 18261 6012
rect 18317 6010 18341 6012
rect 18397 6010 18403 6012
rect 18157 5958 18159 6010
rect 18339 5958 18341 6010
rect 18095 5956 18101 5958
rect 18157 5956 18181 5958
rect 18237 5956 18261 5958
rect 18317 5956 18341 5958
rect 18397 5956 18403 5958
rect 18095 5947 18403 5956
rect 12380 5468 12688 5477
rect 12380 5466 12386 5468
rect 12442 5466 12466 5468
rect 12522 5466 12546 5468
rect 12602 5466 12626 5468
rect 12682 5466 12688 5468
rect 12442 5414 12444 5466
rect 12624 5414 12626 5466
rect 12380 5412 12386 5414
rect 12442 5412 12466 5414
rect 12522 5412 12546 5414
rect 12602 5412 12626 5414
rect 12682 5412 12688 5414
rect 12380 5403 12688 5412
rect 23810 5468 24118 5477
rect 23810 5466 23816 5468
rect 23872 5466 23896 5468
rect 23952 5466 23976 5468
rect 24032 5466 24056 5468
rect 24112 5466 24118 5468
rect 23872 5414 23874 5466
rect 24054 5414 24056 5466
rect 23810 5412 23816 5414
rect 23872 5412 23896 5414
rect 23952 5412 23976 5414
rect 24032 5412 24056 5414
rect 24112 5412 24118 5414
rect 23810 5403 24118 5412
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 6665 4924 6973 4933
rect 6665 4922 6671 4924
rect 6727 4922 6751 4924
rect 6807 4922 6831 4924
rect 6887 4922 6911 4924
rect 6967 4922 6973 4924
rect 6727 4870 6729 4922
rect 6909 4870 6911 4922
rect 6665 4868 6671 4870
rect 6727 4868 6751 4870
rect 6807 4868 6831 4870
rect 6887 4868 6911 4870
rect 6967 4868 6973 4870
rect 6665 4859 6973 4868
rect 18095 4924 18403 4933
rect 18095 4922 18101 4924
rect 18157 4922 18181 4924
rect 18237 4922 18261 4924
rect 18317 4922 18341 4924
rect 18397 4922 18403 4924
rect 18157 4870 18159 4922
rect 18339 4870 18341 4922
rect 18095 4868 18101 4870
rect 18157 4868 18181 4870
rect 18237 4868 18261 4870
rect 18317 4868 18341 4870
rect 18397 4868 18403 4870
rect 18095 4859 18403 4868
rect 12380 4380 12688 4389
rect 12380 4378 12386 4380
rect 12442 4378 12466 4380
rect 12522 4378 12546 4380
rect 12602 4378 12626 4380
rect 12682 4378 12688 4380
rect 12442 4326 12444 4378
rect 12624 4326 12626 4378
rect 12380 4324 12386 4326
rect 12442 4324 12466 4326
rect 12522 4324 12546 4326
rect 12602 4324 12626 4326
rect 12682 4324 12688 4326
rect 12380 4315 12688 4324
rect 23810 4380 24118 4389
rect 23810 4378 23816 4380
rect 23872 4378 23896 4380
rect 23952 4378 23976 4380
rect 24032 4378 24056 4380
rect 24112 4378 24118 4380
rect 23872 4326 23874 4378
rect 24054 4326 24056 4378
rect 23810 4324 23816 4326
rect 23872 4324 23896 4326
rect 23952 4324 23976 4326
rect 24032 4324 24056 4326
rect 24112 4324 24118 4326
rect 23810 4315 24118 4324
rect 6665 3836 6973 3845
rect 6665 3834 6671 3836
rect 6727 3834 6751 3836
rect 6807 3834 6831 3836
rect 6887 3834 6911 3836
rect 6967 3834 6973 3836
rect 6727 3782 6729 3834
rect 6909 3782 6911 3834
rect 6665 3780 6671 3782
rect 6727 3780 6751 3782
rect 6807 3780 6831 3782
rect 6887 3780 6911 3782
rect 6967 3780 6973 3782
rect 6665 3771 6973 3780
rect 18095 3836 18403 3845
rect 18095 3834 18101 3836
rect 18157 3834 18181 3836
rect 18237 3834 18261 3836
rect 18317 3834 18341 3836
rect 18397 3834 18403 3836
rect 18157 3782 18159 3834
rect 18339 3782 18341 3834
rect 18095 3780 18101 3782
rect 18157 3780 18181 3782
rect 18237 3780 18261 3782
rect 18317 3780 18341 3782
rect 18397 3780 18403 3782
rect 18095 3771 18403 3780
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 23664 3596 23716 3602
rect 23664 3538 23716 3544
rect 12380 3292 12688 3301
rect 12380 3290 12386 3292
rect 12442 3290 12466 3292
rect 12522 3290 12546 3292
rect 12602 3290 12626 3292
rect 12682 3290 12688 3292
rect 12442 3238 12444 3290
rect 12624 3238 12626 3290
rect 12380 3236 12386 3238
rect 12442 3236 12466 3238
rect 12522 3236 12546 3238
rect 12602 3236 12626 3238
rect 12682 3236 12688 3238
rect 12380 3227 12688 3236
rect 6665 2748 6973 2757
rect 6665 2746 6671 2748
rect 6727 2746 6751 2748
rect 6807 2746 6831 2748
rect 6887 2746 6911 2748
rect 6967 2746 6973 2748
rect 6727 2694 6729 2746
rect 6909 2694 6911 2746
rect 6665 2692 6671 2694
rect 6727 2692 6751 2694
rect 6807 2692 6831 2694
rect 6887 2692 6911 2694
rect 6967 2692 6973 2694
rect 6665 2683 6973 2692
rect 18095 2748 18403 2757
rect 18095 2746 18101 2748
rect 18157 2746 18181 2748
rect 18237 2746 18261 2748
rect 18317 2746 18341 2748
rect 18397 2746 18403 2748
rect 18157 2694 18159 2746
rect 18339 2694 18341 2746
rect 18095 2692 18101 2694
rect 18157 2692 18181 2694
rect 18237 2692 18261 2694
rect 18317 2692 18341 2694
rect 18397 2692 18403 2694
rect 18095 2683 18403 2692
rect 23676 2650 23704 3538
rect 23810 3292 24118 3301
rect 23810 3290 23816 3292
rect 23872 3290 23896 3292
rect 23952 3290 23976 3292
rect 24032 3290 24056 3292
rect 24112 3290 24118 3292
rect 23872 3238 23874 3290
rect 24054 3238 24056 3290
rect 23810 3236 23816 3238
rect 23872 3236 23896 3238
rect 23952 3236 23976 3238
rect 24032 3236 24056 3238
rect 24112 3236 24118 3238
rect 23810 3227 24118 3236
rect 24228 2650 24256 3606
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 12380 2204 12688 2213
rect 12380 2202 12386 2204
rect 12442 2202 12466 2204
rect 12522 2202 12546 2204
rect 12602 2202 12626 2204
rect 12682 2202 12688 2204
rect 12442 2150 12444 2202
rect 12624 2150 12626 2202
rect 12380 2148 12386 2150
rect 12442 2148 12466 2150
rect 12522 2148 12546 2150
rect 12602 2148 12626 2150
rect 12682 2148 12688 2150
rect 12380 2139 12688 2148
rect 21100 2106 21128 2314
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 21192 2106 21220 2246
rect 22388 2106 22416 2382
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 23216 2106 23244 2314
rect 23492 2106 23520 2518
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 23572 2372 23624 2378
rect 23572 2314 23624 2320
rect 21088 2100 21140 2106
rect 21088 2042 21140 2048
rect 21180 2100 21232 2106
rect 21180 2042 21232 2048
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 23480 2100 23532 2106
rect 23480 2042 23532 2048
rect 20076 1964 20128 1970
rect 20076 1906 20128 1912
rect 20904 1964 20956 1970
rect 20904 1906 20956 1912
rect 22468 1964 22520 1970
rect 22468 1906 22520 1912
rect 22928 1964 22980 1970
rect 22928 1906 22980 1912
rect 23480 1964 23532 1970
rect 23480 1906 23532 1912
rect 19892 1896 19944 1902
rect 19892 1838 19944 1844
rect 6665 1660 6973 1669
rect 6665 1658 6671 1660
rect 6727 1658 6751 1660
rect 6807 1658 6831 1660
rect 6887 1658 6911 1660
rect 6967 1658 6973 1660
rect 6727 1606 6729 1658
rect 6909 1606 6911 1658
rect 6665 1604 6671 1606
rect 6727 1604 6751 1606
rect 6807 1604 6831 1606
rect 6887 1604 6911 1606
rect 6967 1604 6973 1606
rect 6665 1595 6973 1604
rect 18095 1660 18403 1669
rect 18095 1658 18101 1660
rect 18157 1658 18181 1660
rect 18237 1658 18261 1660
rect 18317 1658 18341 1660
rect 18397 1658 18403 1660
rect 18157 1606 18159 1658
rect 18339 1606 18341 1658
rect 18095 1604 18101 1606
rect 18157 1604 18181 1606
rect 18237 1604 18261 1606
rect 18317 1604 18341 1606
rect 18397 1604 18403 1606
rect 18095 1595 18403 1604
rect 15384 1488 15436 1494
rect 15384 1430 15436 1436
rect 1952 1352 2004 1358
rect 1952 1294 2004 1300
rect 4160 1352 4212 1358
rect 4160 1294 4212 1300
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 10784 1352 10836 1358
rect 10784 1294 10836 1300
rect 12992 1352 13044 1358
rect 12992 1294 13044 1300
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 1858 82 1914 160
rect 1964 82 1992 1294
rect 2136 1216 2188 1222
rect 2136 1158 2188 1164
rect 2148 1018 2176 1158
rect 2136 1012 2188 1018
rect 2136 954 2188 960
rect 1858 54 1992 82
rect 4066 82 4122 160
rect 4172 82 4200 1294
rect 4066 54 4200 82
rect 6274 82 6330 160
rect 6380 82 6408 1294
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 6564 950 6592 1158
rect 6552 944 6604 950
rect 6552 886 6604 892
rect 6274 54 6408 82
rect 8482 82 8538 160
rect 8588 82 8616 1294
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8772 1018 8800 1158
rect 8760 1012 8812 1018
rect 8760 954 8812 960
rect 8482 54 8616 82
rect 10690 82 10746 160
rect 10796 82 10824 1294
rect 10968 1216 11020 1222
rect 10968 1158 11020 1164
rect 10980 746 11008 1158
rect 12380 1116 12688 1125
rect 12380 1114 12386 1116
rect 12442 1114 12466 1116
rect 12522 1114 12546 1116
rect 12602 1114 12626 1116
rect 12682 1114 12688 1116
rect 12442 1062 12444 1114
rect 12624 1062 12626 1114
rect 12380 1060 12386 1062
rect 12442 1060 12466 1062
rect 12522 1060 12546 1062
rect 12602 1060 12626 1062
rect 12682 1060 12688 1062
rect 12380 1051 12688 1060
rect 10968 740 11020 746
rect 10968 682 11020 688
rect 10690 54 10824 82
rect 12898 82 12954 160
rect 13004 82 13032 1294
rect 12898 54 13032 82
rect 15106 82 15162 160
rect 15212 82 15240 1294
rect 15396 950 15424 1430
rect 17408 1352 17460 1358
rect 17408 1294 17460 1300
rect 19616 1352 19668 1358
rect 19616 1294 19668 1300
rect 15476 1216 15528 1222
rect 15476 1158 15528 1164
rect 15488 950 15516 1158
rect 15384 944 15436 950
rect 15384 886 15436 892
rect 15476 944 15528 950
rect 15476 886 15528 892
rect 15106 54 15240 82
rect 17314 82 17370 160
rect 17420 82 17448 1294
rect 17314 54 17448 82
rect 19522 82 19578 160
rect 19628 82 19656 1294
rect 19904 1018 19932 1838
rect 20088 1562 20116 1906
rect 20076 1556 20128 1562
rect 20076 1498 20128 1504
rect 20916 1290 20944 1906
rect 22480 1562 22508 1906
rect 22468 1556 22520 1562
rect 22468 1498 22520 1504
rect 21824 1352 21876 1358
rect 21824 1294 21876 1300
rect 20904 1284 20956 1290
rect 20904 1226 20956 1232
rect 21180 1284 21232 1290
rect 21180 1226 21232 1232
rect 21192 1018 21220 1226
rect 19892 1012 19944 1018
rect 19892 954 19944 960
rect 21180 1012 21232 1018
rect 21180 954 21232 960
rect 19522 54 19656 82
rect 21730 82 21786 160
rect 21836 82 21864 1294
rect 22940 678 22968 1906
rect 23296 1896 23348 1902
rect 23296 1838 23348 1844
rect 23204 1352 23256 1358
rect 23204 1294 23256 1300
rect 23216 1018 23244 1294
rect 23204 1012 23256 1018
rect 23204 954 23256 960
rect 23308 746 23336 1838
rect 23492 1222 23520 1906
rect 23584 1562 23612 2314
rect 23676 1850 23704 2382
rect 23810 2204 24118 2213
rect 23810 2202 23816 2204
rect 23872 2202 23896 2204
rect 23952 2202 23976 2204
rect 24032 2202 24056 2204
rect 24112 2202 24118 2204
rect 23872 2150 23874 2202
rect 24054 2150 24056 2202
rect 23810 2148 23816 2150
rect 23872 2148 23896 2150
rect 23952 2148 23976 2150
rect 24032 2148 24056 2150
rect 24112 2148 24118 2150
rect 23810 2139 24118 2148
rect 24596 2106 24624 2382
rect 24584 2100 24636 2106
rect 24584 2042 24636 2048
rect 24032 1964 24084 1970
rect 24032 1906 24084 1912
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 23676 1834 23796 1850
rect 23676 1828 23808 1834
rect 23676 1822 23756 1828
rect 23756 1770 23808 1776
rect 24044 1562 24072 1906
rect 24504 1562 24532 1906
rect 24688 1766 24716 4966
rect 24780 2650 24808 6122
rect 29525 6012 29833 6021
rect 29525 6010 29531 6012
rect 29587 6010 29611 6012
rect 29667 6010 29691 6012
rect 29747 6010 29771 6012
rect 29827 6010 29833 6012
rect 29587 5958 29589 6010
rect 29769 5958 29771 6010
rect 29525 5956 29531 5958
rect 29587 5956 29611 5958
rect 29667 5956 29691 5958
rect 29747 5956 29771 5958
rect 29827 5956 29833 5958
rect 29525 5947 29833 5956
rect 32128 5636 32180 5642
rect 32128 5578 32180 5584
rect 29525 4924 29833 4933
rect 29525 4922 29531 4924
rect 29587 4922 29611 4924
rect 29667 4922 29691 4924
rect 29747 4922 29771 4924
rect 29827 4922 29833 4924
rect 29587 4870 29589 4922
rect 29769 4870 29771 4922
rect 29525 4868 29531 4870
rect 29587 4868 29611 4870
rect 29667 4868 29691 4870
rect 29747 4868 29771 4870
rect 29827 4868 29833 4870
rect 29525 4859 29833 4868
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 25688 3460 25740 3466
rect 25688 3402 25740 3408
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24780 2514 24992 2530
rect 24768 2508 24992 2514
rect 24820 2502 24992 2508
rect 24768 2450 24820 2456
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24872 1970 24900 2382
rect 24964 2310 24992 2502
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 25424 2106 25452 2382
rect 25412 2100 25464 2106
rect 25412 2042 25464 2048
rect 24768 1964 24820 1970
rect 24768 1906 24820 1912
rect 24860 1964 24912 1970
rect 24860 1906 24912 1912
rect 24676 1760 24728 1766
rect 24676 1702 24728 1708
rect 23572 1556 23624 1562
rect 23572 1498 23624 1504
rect 24032 1556 24084 1562
rect 24032 1498 24084 1504
rect 24492 1556 24544 1562
rect 24492 1498 24544 1504
rect 24032 1352 24084 1358
rect 24084 1312 24256 1340
rect 24032 1294 24084 1300
rect 23480 1216 23532 1222
rect 23480 1158 23532 1164
rect 23810 1116 24118 1125
rect 23810 1114 23816 1116
rect 23872 1114 23896 1116
rect 23952 1114 23976 1116
rect 24032 1114 24056 1116
rect 24112 1114 24118 1116
rect 23872 1062 23874 1114
rect 24054 1062 24056 1114
rect 23810 1060 23816 1062
rect 23872 1060 23896 1062
rect 23952 1060 23976 1062
rect 24032 1060 24056 1062
rect 24112 1060 24118 1062
rect 23810 1051 24118 1060
rect 23296 740 23348 746
rect 23296 682 23348 688
rect 22928 672 22980 678
rect 22928 614 22980 620
rect 21730 54 21864 82
rect 23938 82 23994 160
rect 24228 82 24256 1312
rect 24780 814 24808 1906
rect 25700 1834 25728 3402
rect 27724 2650 27752 4762
rect 29525 3836 29833 3845
rect 29525 3834 29531 3836
rect 29587 3834 29611 3836
rect 29667 3834 29691 3836
rect 29747 3834 29771 3836
rect 29827 3834 29833 3836
rect 29587 3782 29589 3834
rect 29769 3782 29771 3834
rect 29525 3780 29531 3782
rect 29587 3780 29611 3782
rect 29667 3780 29691 3782
rect 29747 3780 29771 3782
rect 29827 3780 29833 3782
rect 29525 3771 29833 3780
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29525 2748 29833 2757
rect 29525 2746 29531 2748
rect 29587 2746 29611 2748
rect 29667 2746 29691 2748
rect 29747 2746 29771 2748
rect 29827 2746 29833 2748
rect 29587 2694 29589 2746
rect 29769 2694 29771 2746
rect 29525 2692 29531 2694
rect 29587 2692 29611 2694
rect 29667 2692 29691 2694
rect 29747 2692 29771 2694
rect 29827 2692 29833 2694
rect 29525 2683 29833 2692
rect 29932 2650 29960 3470
rect 32140 2650 32168 5578
rect 33704 3670 33732 8366
rect 33692 3664 33744 3670
rect 33692 3606 33744 3612
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 27712 2644 27764 2650
rect 27712 2586 27764 2592
rect 29920 2644 29972 2650
rect 29920 2586 29972 2592
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 27540 2106 27568 2382
rect 27528 2100 27580 2106
rect 27528 2042 27580 2048
rect 26976 1964 27028 1970
rect 26976 1906 27028 1912
rect 25688 1828 25740 1834
rect 25688 1770 25740 1776
rect 26988 1562 27016 1906
rect 27632 1766 27660 2586
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 29748 2106 29776 2382
rect 31404 2106 31432 2382
rect 33888 2310 33916 9318
rect 34060 9308 34112 9314
rect 34060 9250 34112 9256
rect 33968 9172 34020 9178
rect 33968 9114 34020 9120
rect 33980 8634 34008 9114
rect 34072 8634 34100 9250
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 34164 8498 34192 9846
rect 34242 9840 34298 10000
rect 34610 9840 34666 10000
rect 34716 9846 34928 9874
rect 34716 9840 34744 9846
rect 34256 8498 34284 9840
rect 34624 9812 34744 9840
rect 34336 9716 34388 9722
rect 34336 9658 34388 9664
rect 34348 9178 34376 9658
rect 34612 9308 34664 9314
rect 34612 9250 34664 9256
rect 34336 9172 34388 9178
rect 34336 9114 34388 9120
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34244 8492 34296 8498
rect 34244 8434 34296 8440
rect 34532 6186 34560 8774
rect 34520 6180 34572 6186
rect 34520 6122 34572 6128
rect 34624 5030 34652 9250
rect 34900 8498 34928 9846
rect 34978 9840 35034 10000
rect 35072 9988 35124 9994
rect 35072 9930 35124 9936
rect 34992 8498 35020 9840
rect 35084 8634 35112 9930
rect 35346 9840 35402 10000
rect 35452 9846 35664 9874
rect 35452 9840 35480 9846
rect 35360 9812 35480 9840
rect 35240 8732 35548 8741
rect 35240 8730 35246 8732
rect 35302 8730 35326 8732
rect 35382 8730 35406 8732
rect 35462 8730 35486 8732
rect 35542 8730 35548 8732
rect 35302 8678 35304 8730
rect 35484 8678 35486 8730
rect 35240 8676 35246 8678
rect 35302 8676 35326 8678
rect 35382 8676 35406 8678
rect 35462 8676 35486 8678
rect 35542 8676 35548 8678
rect 35240 8667 35548 8676
rect 35072 8628 35124 8634
rect 35072 8570 35124 8576
rect 35636 8498 35664 9846
rect 35714 9840 35770 10000
rect 36082 9840 36138 10000
rect 36188 9846 36400 9874
rect 36188 9840 36216 9846
rect 35728 8498 35756 9840
rect 36096 9812 36216 9840
rect 36176 8900 36228 8906
rect 36176 8842 36228 8848
rect 36268 8900 36320 8906
rect 36268 8842 36320 8848
rect 36188 8634 36216 8842
rect 36176 8628 36228 8634
rect 36176 8570 36228 8576
rect 34888 8492 34940 8498
rect 34888 8434 34940 8440
rect 34980 8492 35032 8498
rect 34980 8434 35032 8440
rect 35624 8492 35676 8498
rect 35624 8434 35676 8440
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35072 8356 35124 8362
rect 35072 8298 35124 8304
rect 35808 8356 35860 8362
rect 35808 8298 35860 8304
rect 35084 8129 35112 8298
rect 35070 8120 35126 8129
rect 35070 8055 35126 8064
rect 35820 7993 35848 8298
rect 35806 7984 35862 7993
rect 35806 7919 35862 7928
rect 35240 7644 35548 7653
rect 35240 7642 35246 7644
rect 35302 7642 35326 7644
rect 35382 7642 35406 7644
rect 35462 7642 35486 7644
rect 35542 7642 35548 7644
rect 35302 7590 35304 7642
rect 35484 7590 35486 7642
rect 35240 7588 35246 7590
rect 35302 7588 35326 7590
rect 35382 7588 35406 7590
rect 35462 7588 35486 7590
rect 35542 7588 35548 7590
rect 35240 7579 35548 7588
rect 36280 6914 36308 8842
rect 36372 8498 36400 9846
rect 36450 9840 36506 10000
rect 36556 9846 36768 9874
rect 36556 9840 36584 9846
rect 36464 9812 36584 9840
rect 36452 9172 36504 9178
rect 36452 9114 36504 9120
rect 36360 8492 36412 8498
rect 36360 8434 36412 8440
rect 36464 8362 36492 9114
rect 36636 9104 36688 9110
rect 36636 9046 36688 9052
rect 36544 9036 36596 9042
rect 36544 8978 36596 8984
rect 36556 8634 36584 8978
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 36452 8356 36504 8362
rect 36452 8298 36504 8304
rect 36452 7336 36504 7342
rect 36452 7278 36504 7284
rect 36096 6886 36308 6914
rect 35240 6556 35548 6565
rect 35240 6554 35246 6556
rect 35302 6554 35326 6556
rect 35382 6554 35406 6556
rect 35462 6554 35486 6556
rect 35542 6554 35548 6556
rect 35302 6502 35304 6554
rect 35484 6502 35486 6554
rect 35240 6500 35246 6502
rect 35302 6500 35326 6502
rect 35382 6500 35406 6502
rect 35462 6500 35486 6502
rect 35542 6500 35548 6502
rect 35240 6491 35548 6500
rect 35240 5468 35548 5477
rect 35240 5466 35246 5468
rect 35302 5466 35326 5468
rect 35382 5466 35406 5468
rect 35462 5466 35486 5468
rect 35542 5466 35548 5468
rect 35302 5414 35304 5466
rect 35484 5414 35486 5466
rect 35240 5412 35246 5414
rect 35302 5412 35326 5414
rect 35382 5412 35406 5414
rect 35462 5412 35486 5414
rect 35542 5412 35548 5414
rect 35240 5403 35548 5412
rect 34612 5024 34664 5030
rect 34612 4966 34664 4972
rect 35240 4380 35548 4389
rect 35240 4378 35246 4380
rect 35302 4378 35326 4380
rect 35382 4378 35406 4380
rect 35462 4378 35486 4380
rect 35542 4378 35548 4380
rect 35302 4326 35304 4378
rect 35484 4326 35486 4378
rect 35240 4324 35246 4326
rect 35302 4324 35326 4326
rect 35382 4324 35406 4326
rect 35462 4324 35486 4326
rect 35542 4324 35548 4326
rect 35240 4315 35548 4324
rect 36096 3602 36124 6886
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 35240 3292 35548 3301
rect 35240 3290 35246 3292
rect 35302 3290 35326 3292
rect 35382 3290 35406 3292
rect 35462 3290 35486 3292
rect 35542 3290 35548 3292
rect 35302 3238 35304 3290
rect 35484 3238 35486 3290
rect 35240 3236 35246 3238
rect 35302 3236 35326 3238
rect 35382 3236 35406 3238
rect 35462 3236 35486 3238
rect 35542 3236 35548 3238
rect 35240 3227 35548 3236
rect 36464 2650 36492 7278
rect 36648 5642 36676 9046
rect 36740 8498 36768 9846
rect 36818 9840 36874 10000
rect 36924 9846 37136 9874
rect 36924 9840 36952 9846
rect 36832 9812 36952 9840
rect 36820 9036 36872 9042
rect 36820 8978 36872 8984
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36636 5636 36688 5642
rect 36636 5578 36688 5584
rect 36452 2644 36504 2650
rect 36452 2586 36504 2592
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 36452 2440 36504 2446
rect 36452 2382 36504 2388
rect 33876 2304 33928 2310
rect 33876 2246 33928 2252
rect 34164 2106 34192 2382
rect 35240 2204 35548 2213
rect 35240 2202 35246 2204
rect 35302 2202 35326 2204
rect 35382 2202 35406 2204
rect 35462 2202 35486 2204
rect 35542 2202 35548 2204
rect 35302 2150 35304 2202
rect 35484 2150 35486 2202
rect 35240 2148 35246 2150
rect 35302 2148 35326 2150
rect 35382 2148 35406 2150
rect 35462 2148 35486 2150
rect 35542 2148 35548 2150
rect 35240 2139 35548 2148
rect 36464 2106 36492 2382
rect 29736 2100 29788 2106
rect 29736 2042 29788 2048
rect 31392 2100 31444 2106
rect 31392 2042 31444 2048
rect 34152 2100 34204 2106
rect 34152 2042 34204 2048
rect 36452 2100 36504 2106
rect 36452 2042 36504 2048
rect 29092 1964 29144 1970
rect 29092 1906 29144 1912
rect 31208 1964 31260 1970
rect 31208 1906 31260 1912
rect 33508 1964 33560 1970
rect 33508 1906 33560 1912
rect 35532 1964 35584 1970
rect 35532 1906 35584 1912
rect 27620 1760 27672 1766
rect 27620 1702 27672 1708
rect 29104 1562 29132 1906
rect 29525 1660 29833 1669
rect 29525 1658 29531 1660
rect 29587 1658 29611 1660
rect 29667 1658 29691 1660
rect 29747 1658 29771 1660
rect 29827 1658 29833 1660
rect 29587 1606 29589 1658
rect 29769 1606 29771 1658
rect 29525 1604 29531 1606
rect 29587 1604 29611 1606
rect 29667 1604 29691 1606
rect 29747 1604 29771 1606
rect 29827 1604 29833 1606
rect 29525 1595 29833 1604
rect 31220 1562 31248 1906
rect 33520 1562 33548 1906
rect 35544 1562 35572 1906
rect 36832 1766 36860 8978
rect 37004 8968 37056 8974
rect 37004 8910 37056 8916
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 36924 7274 36952 8570
rect 37016 8362 37044 8910
rect 37108 8498 37136 9846
rect 37186 9840 37242 10000
rect 37554 9840 37610 10000
rect 37660 9846 37872 9874
rect 37660 9840 37688 9846
rect 37200 8498 37228 9840
rect 37568 9812 37688 9840
rect 37648 9648 37700 9654
rect 37648 9590 37700 9596
rect 37096 8492 37148 8498
rect 37096 8434 37148 8440
rect 37188 8492 37240 8498
rect 37188 8434 37240 8440
rect 37004 8356 37056 8362
rect 37004 8298 37056 8304
rect 37096 8356 37148 8362
rect 37096 8298 37148 8304
rect 37108 7818 37136 8298
rect 37660 8294 37688 9590
rect 37844 8498 37872 9846
rect 37922 9840 37978 10000
rect 38028 9846 38240 9874
rect 38028 9840 38056 9846
rect 37936 9812 38056 9840
rect 38212 8498 38240 9846
rect 38290 9840 38346 10000
rect 38396 9846 38608 9874
rect 38396 9840 38424 9846
rect 38304 9812 38424 9840
rect 38580 8498 38608 9846
rect 38658 9840 38714 10000
rect 38764 9846 38976 9874
rect 38764 9840 38792 9846
rect 38672 9812 38792 9840
rect 38948 8498 38976 9846
rect 39026 9840 39082 10000
rect 39132 9846 39344 9874
rect 39132 9840 39160 9846
rect 39040 9812 39160 9840
rect 39120 9240 39172 9246
rect 39120 9182 39172 9188
rect 39132 8634 39160 9182
rect 39120 8628 39172 8634
rect 39120 8570 39172 8576
rect 39316 8498 39344 9846
rect 39394 9840 39450 10000
rect 39762 9840 39818 10000
rect 40130 9840 40186 10000
rect 40498 9840 40554 10000
rect 40866 9840 40922 10000
rect 41234 9840 41290 10000
rect 41602 9840 41658 10000
rect 41970 9840 42026 10000
rect 42338 9840 42394 10000
rect 42444 9846 42656 9874
rect 42444 9840 42472 9846
rect 39408 8634 39436 9840
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 39776 8566 39804 9840
rect 39764 8560 39816 8566
rect 39764 8502 39816 8508
rect 37832 8492 37884 8498
rect 37832 8434 37884 8440
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 38568 8492 38620 8498
rect 38568 8434 38620 8440
rect 38936 8492 38988 8498
rect 38936 8434 38988 8440
rect 39304 8492 39356 8498
rect 39304 8434 39356 8440
rect 39948 8492 40000 8498
rect 39948 8434 40000 8440
rect 38752 8356 38804 8362
rect 38752 8298 38804 8304
rect 37648 8288 37700 8294
rect 37648 8230 37700 8236
rect 37096 7812 37148 7818
rect 37096 7754 37148 7760
rect 38764 7449 38792 8298
rect 38750 7440 38806 7449
rect 38750 7375 38806 7384
rect 36912 7268 36964 7274
rect 36912 7210 36964 7216
rect 39960 3466 39988 8434
rect 40144 8362 40172 9840
rect 40224 8492 40276 8498
rect 40224 8434 40276 8440
rect 40132 8356 40184 8362
rect 40132 8298 40184 8304
rect 40040 7880 40092 7886
rect 40040 7822 40092 7828
rect 39948 3460 40000 3466
rect 39948 3402 40000 3408
rect 40052 2514 40080 7822
rect 40236 2514 40264 8434
rect 40512 8090 40540 9840
rect 40684 8832 40736 8838
rect 40684 8774 40736 8780
rect 40696 8634 40724 8774
rect 40880 8634 40908 9840
rect 40684 8628 40736 8634
rect 40684 8570 40736 8576
rect 40868 8628 40920 8634
rect 40868 8570 40920 8576
rect 41248 8566 41276 9840
rect 41236 8560 41288 8566
rect 41236 8502 41288 8508
rect 40592 8492 40644 8498
rect 40592 8434 40644 8440
rect 40500 8084 40552 8090
rect 40500 8026 40552 8032
rect 40040 2508 40092 2514
rect 40040 2450 40092 2456
rect 40224 2508 40276 2514
rect 40224 2450 40276 2456
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38672 2106 38700 2382
rect 40604 2378 40632 8434
rect 41616 8362 41644 9840
rect 41984 8430 42012 9840
rect 42352 9812 42472 9840
rect 41972 8424 42024 8430
rect 41972 8366 42024 8372
rect 41604 8356 41656 8362
rect 41604 8298 41656 8304
rect 42628 8242 42656 9846
rect 42706 9840 42762 10000
rect 43074 9840 43130 10000
rect 43180 9846 43392 9874
rect 43180 9840 43208 9846
rect 42720 8634 42748 9840
rect 43088 9812 43208 9840
rect 42800 9308 42852 9314
rect 42800 9250 42852 9256
rect 42708 8628 42760 8634
rect 42708 8570 42760 8576
rect 42812 8566 42840 9250
rect 43364 8566 43392 9846
rect 43442 9840 43498 10000
rect 43548 9846 43760 9874
rect 43548 9840 43576 9846
rect 43456 9812 43576 9840
rect 43628 8900 43680 8906
rect 43628 8842 43680 8848
rect 42800 8560 42852 8566
rect 42800 8502 42852 8508
rect 43352 8560 43404 8566
rect 43352 8502 43404 8508
rect 43640 8498 43668 8842
rect 43628 8492 43680 8498
rect 43628 8434 43680 8440
rect 42628 8214 42840 8242
rect 40955 8188 41263 8197
rect 40955 8186 40961 8188
rect 41017 8186 41041 8188
rect 41097 8186 41121 8188
rect 41177 8186 41201 8188
rect 41257 8186 41263 8188
rect 41017 8134 41019 8186
rect 41199 8134 41201 8186
rect 40955 8132 40961 8134
rect 41017 8132 41041 8134
rect 41097 8132 41121 8134
rect 41177 8132 41201 8134
rect 41257 8132 41263 8134
rect 40955 8123 41263 8132
rect 42812 8090 42840 8214
rect 43732 8090 43760 9846
rect 43810 9840 43866 10000
rect 43916 9846 44128 9874
rect 43916 9840 43944 9846
rect 43824 9812 43944 9840
rect 43812 9376 43864 9382
rect 43812 9318 43864 9324
rect 43824 8498 43852 9318
rect 43812 8492 43864 8498
rect 43812 8434 43864 8440
rect 44100 8242 44128 9846
rect 44178 9840 44234 10000
rect 44284 9846 44496 9874
rect 44284 9840 44312 9846
rect 44192 9812 44312 9840
rect 44468 8634 44496 9846
rect 44546 9840 44602 10000
rect 44914 9840 44970 10000
rect 45282 9840 45338 10000
rect 45650 9840 45706 10000
rect 46018 9840 46074 10000
rect 46386 9840 46442 10000
rect 46754 9840 46810 10000
rect 44456 8628 44508 8634
rect 44456 8570 44508 8576
rect 44100 8214 44220 8242
rect 42800 8084 42852 8090
rect 42800 8026 42852 8032
rect 43720 8084 43772 8090
rect 43720 8026 43772 8032
rect 44192 8022 44220 8214
rect 44180 8016 44232 8022
rect 44180 7958 44232 7964
rect 43260 7812 43312 7818
rect 43260 7754 43312 7760
rect 43996 7812 44048 7818
rect 43996 7754 44048 7760
rect 41604 7404 41656 7410
rect 41604 7346 41656 7352
rect 40955 7100 41263 7109
rect 40955 7098 40961 7100
rect 41017 7098 41041 7100
rect 41097 7098 41121 7100
rect 41177 7098 41201 7100
rect 41257 7098 41263 7100
rect 41017 7046 41019 7098
rect 41199 7046 41201 7098
rect 40955 7044 40961 7046
rect 41017 7044 41041 7046
rect 41097 7044 41121 7046
rect 41177 7044 41201 7046
rect 41257 7044 41263 7046
rect 40955 7035 41263 7044
rect 40955 6012 41263 6021
rect 40955 6010 40961 6012
rect 41017 6010 41041 6012
rect 41097 6010 41121 6012
rect 41177 6010 41201 6012
rect 41257 6010 41263 6012
rect 41017 5958 41019 6010
rect 41199 5958 41201 6010
rect 40955 5956 40961 5958
rect 41017 5956 41041 5958
rect 41097 5956 41121 5958
rect 41177 5956 41201 5958
rect 41257 5956 41263 5958
rect 40955 5947 41263 5956
rect 40955 4924 41263 4933
rect 40955 4922 40961 4924
rect 41017 4922 41041 4924
rect 41097 4922 41121 4924
rect 41177 4922 41201 4924
rect 41257 4922 41263 4924
rect 41017 4870 41019 4922
rect 41199 4870 41201 4922
rect 40955 4868 40961 4870
rect 41017 4868 41041 4870
rect 41097 4868 41121 4870
rect 41177 4868 41201 4870
rect 41257 4868 41263 4870
rect 40955 4859 41263 4868
rect 40955 3836 41263 3845
rect 40955 3834 40961 3836
rect 41017 3834 41041 3836
rect 41097 3834 41121 3836
rect 41177 3834 41201 3836
rect 41257 3834 41263 3836
rect 41017 3782 41019 3834
rect 41199 3782 41201 3834
rect 40955 3780 40961 3782
rect 41017 3780 41041 3782
rect 41097 3780 41121 3782
rect 41177 3780 41201 3782
rect 41257 3780 41263 3782
rect 40955 3771 41263 3780
rect 40955 2748 41263 2757
rect 40955 2746 40961 2748
rect 41017 2746 41041 2748
rect 41097 2746 41121 2748
rect 41177 2746 41201 2748
rect 41257 2746 41263 2748
rect 41017 2694 41019 2746
rect 41199 2694 41201 2746
rect 40955 2692 40961 2694
rect 41017 2692 41041 2694
rect 41097 2692 41121 2694
rect 41177 2692 41201 2694
rect 41257 2692 41263 2694
rect 40955 2683 41263 2692
rect 41616 2650 41644 7346
rect 42800 6724 42852 6730
rect 42800 6666 42852 6672
rect 42812 2650 42840 6666
rect 41604 2644 41656 2650
rect 41604 2586 41656 2592
rect 42800 2644 42852 2650
rect 42800 2586 42852 2592
rect 43076 2440 43128 2446
rect 43076 2382 43128 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 43088 2106 43116 2382
rect 43272 2106 43300 7754
rect 44008 3534 44036 7754
rect 44560 7546 44588 9840
rect 44548 7540 44600 7546
rect 44548 7482 44600 7488
rect 44928 6866 44956 9840
rect 45100 9036 45152 9042
rect 45100 8978 45152 8984
rect 45112 8498 45140 8978
rect 45100 8492 45152 8498
rect 45100 8434 45152 8440
rect 45100 7812 45152 7818
rect 45100 7754 45152 7760
rect 44916 6860 44968 6866
rect 44916 6802 44968 6808
rect 44364 6792 44416 6798
rect 44364 6734 44416 6740
rect 43996 3528 44048 3534
rect 43996 3470 44048 3476
rect 44376 2650 44404 6734
rect 45112 4826 45140 7754
rect 45296 7546 45324 9840
rect 45468 9104 45520 9110
rect 45468 9046 45520 9052
rect 45480 8566 45508 9046
rect 45468 8560 45520 8566
rect 45468 8502 45520 8508
rect 45664 7546 45692 9840
rect 45836 7812 45888 7818
rect 45836 7754 45888 7760
rect 45284 7540 45336 7546
rect 45284 7482 45336 7488
rect 45652 7540 45704 7546
rect 45652 7482 45704 7488
rect 45560 7404 45612 7410
rect 45560 7346 45612 7352
rect 45652 7404 45704 7410
rect 45652 7346 45704 7352
rect 45100 4820 45152 4826
rect 45100 4762 45152 4768
rect 45572 2650 45600 7346
rect 45664 2650 45692 7346
rect 45848 6914 45876 7754
rect 46032 7002 46060 9840
rect 46400 7546 46428 9840
rect 46768 8922 46796 9840
rect 46584 8894 46796 8922
rect 46584 8090 46612 8894
rect 46670 8732 46978 8741
rect 46670 8730 46676 8732
rect 46732 8730 46756 8732
rect 46812 8730 46836 8732
rect 46892 8730 46916 8732
rect 46972 8730 46978 8732
rect 46732 8678 46734 8730
rect 46914 8678 46916 8730
rect 46670 8676 46676 8678
rect 46732 8676 46756 8678
rect 46812 8676 46836 8678
rect 46892 8676 46916 8678
rect 46972 8676 46978 8678
rect 46670 8667 46978 8676
rect 46572 8084 46624 8090
rect 46572 8026 46624 8032
rect 46670 7644 46978 7653
rect 46670 7642 46676 7644
rect 46732 7642 46756 7644
rect 46812 7642 46836 7644
rect 46892 7642 46916 7644
rect 46972 7642 46978 7644
rect 46732 7590 46734 7642
rect 46914 7590 46916 7642
rect 46670 7588 46676 7590
rect 46732 7588 46756 7590
rect 46812 7588 46836 7590
rect 46892 7588 46916 7590
rect 46972 7588 46978 7590
rect 46670 7579 46978 7588
rect 46388 7540 46440 7546
rect 46388 7482 46440 7488
rect 46020 6996 46072 7002
rect 46020 6938 46072 6944
rect 45756 6886 45876 6914
rect 45756 2650 45784 6886
rect 46670 6556 46978 6565
rect 46670 6554 46676 6556
rect 46732 6554 46756 6556
rect 46812 6554 46836 6556
rect 46892 6554 46916 6556
rect 46972 6554 46978 6556
rect 46732 6502 46734 6554
rect 46914 6502 46916 6554
rect 46670 6500 46676 6502
rect 46732 6500 46756 6502
rect 46812 6500 46836 6502
rect 46892 6500 46916 6502
rect 46972 6500 46978 6502
rect 46670 6491 46978 6500
rect 46670 5468 46978 5477
rect 46670 5466 46676 5468
rect 46732 5466 46756 5468
rect 46812 5466 46836 5468
rect 46892 5466 46916 5468
rect 46972 5466 46978 5468
rect 46732 5414 46734 5466
rect 46914 5414 46916 5466
rect 46670 5412 46676 5414
rect 46732 5412 46756 5414
rect 46812 5412 46836 5414
rect 46892 5412 46916 5414
rect 46972 5412 46978 5414
rect 46670 5403 46978 5412
rect 46670 4380 46978 4389
rect 46670 4378 46676 4380
rect 46732 4378 46756 4380
rect 46812 4378 46836 4380
rect 46892 4378 46916 4380
rect 46972 4378 46978 4380
rect 46732 4326 46734 4378
rect 46914 4326 46916 4378
rect 46670 4324 46676 4326
rect 46732 4324 46756 4326
rect 46812 4324 46836 4326
rect 46892 4324 46916 4326
rect 46972 4324 46978 4326
rect 46670 4315 46978 4324
rect 46670 3292 46978 3301
rect 46670 3290 46676 3292
rect 46732 3290 46756 3292
rect 46812 3290 46836 3292
rect 46892 3290 46916 3292
rect 46972 3290 46978 3292
rect 46732 3238 46734 3290
rect 46914 3238 46916 3290
rect 46670 3236 46676 3238
rect 46732 3236 46756 3238
rect 46812 3236 46836 3238
rect 46892 3236 46916 3238
rect 46972 3236 46978 3238
rect 46670 3227 46978 3236
rect 44364 2644 44416 2650
rect 44364 2586 44416 2592
rect 45560 2644 45612 2650
rect 45560 2586 45612 2592
rect 45652 2644 45704 2650
rect 45652 2586 45704 2592
rect 45744 2644 45796 2650
rect 45744 2586 45796 2592
rect 45008 2440 45060 2446
rect 45008 2382 45060 2388
rect 45928 2440 45980 2446
rect 45928 2382 45980 2388
rect 44732 2372 44784 2378
rect 44732 2314 44784 2320
rect 38660 2100 38712 2106
rect 38660 2042 38712 2048
rect 43076 2100 43128 2106
rect 43076 2042 43128 2048
rect 43260 2100 43312 2106
rect 43260 2042 43312 2048
rect 37740 1964 37792 1970
rect 37740 1906 37792 1912
rect 42432 1964 42484 1970
rect 42432 1906 42484 1912
rect 44088 1964 44140 1970
rect 44088 1906 44140 1912
rect 44548 1964 44600 1970
rect 44548 1906 44600 1912
rect 36820 1760 36872 1766
rect 36820 1702 36872 1708
rect 37752 1562 37780 1906
rect 40955 1660 41263 1669
rect 40955 1658 40961 1660
rect 41017 1658 41041 1660
rect 41097 1658 41121 1660
rect 41177 1658 41201 1660
rect 41257 1658 41263 1660
rect 41017 1606 41019 1658
rect 41199 1606 41201 1658
rect 40955 1604 40961 1606
rect 41017 1604 41041 1606
rect 41097 1604 41121 1606
rect 41177 1604 41201 1606
rect 41257 1604 41263 1606
rect 40955 1595 41263 1604
rect 42444 1562 42472 1906
rect 26976 1556 27028 1562
rect 26976 1498 27028 1504
rect 29092 1556 29144 1562
rect 29092 1498 29144 1504
rect 31208 1556 31260 1562
rect 31208 1498 31260 1504
rect 33508 1556 33560 1562
rect 33508 1498 33560 1504
rect 35532 1556 35584 1562
rect 35532 1498 35584 1504
rect 37740 1556 37792 1562
rect 37740 1498 37792 1504
rect 42432 1556 42484 1562
rect 42432 1498 42484 1504
rect 26240 1352 26292 1358
rect 26240 1294 26292 1300
rect 28448 1352 28500 1358
rect 28448 1294 28500 1300
rect 30656 1352 30708 1358
rect 30656 1294 30708 1300
rect 32864 1352 32916 1358
rect 32864 1294 32916 1300
rect 35072 1352 35124 1358
rect 35072 1294 35124 1300
rect 37280 1352 37332 1358
rect 37280 1294 37332 1300
rect 39488 1352 39540 1358
rect 39488 1294 39540 1300
rect 41696 1352 41748 1358
rect 41696 1294 41748 1300
rect 43904 1352 43956 1358
rect 43904 1294 43956 1300
rect 24768 808 24820 814
rect 26252 762 26280 1294
rect 24768 750 24820 756
rect 26160 734 26280 762
rect 26160 160 26188 734
rect 23938 54 24256 82
rect 1858 0 1914 54
rect 4066 0 4122 54
rect 6274 0 6330 54
rect 8482 0 8538 54
rect 10690 0 10746 54
rect 12898 0 12954 54
rect 15106 0 15162 54
rect 17314 0 17370 54
rect 19522 0 19578 54
rect 21730 0 21786 54
rect 23938 0 23994 54
rect 26146 0 26202 160
rect 28354 82 28410 160
rect 28460 82 28488 1294
rect 28354 54 28488 82
rect 30562 82 30618 160
rect 30668 82 30696 1294
rect 30562 54 30696 82
rect 32770 82 32826 160
rect 32876 82 32904 1294
rect 32770 54 32904 82
rect 34978 82 35034 160
rect 35084 82 35112 1294
rect 35240 1116 35548 1125
rect 35240 1114 35246 1116
rect 35302 1114 35326 1116
rect 35382 1114 35406 1116
rect 35462 1114 35486 1116
rect 35542 1114 35548 1116
rect 35302 1062 35304 1114
rect 35484 1062 35486 1114
rect 35240 1060 35246 1062
rect 35302 1060 35326 1062
rect 35382 1060 35406 1062
rect 35462 1060 35486 1062
rect 35542 1060 35548 1062
rect 35240 1051 35548 1060
rect 34978 54 35112 82
rect 37186 82 37242 160
rect 37292 82 37320 1294
rect 37186 54 37320 82
rect 39394 82 39450 160
rect 39500 82 39528 1294
rect 39394 54 39528 82
rect 41602 82 41658 160
rect 41708 82 41736 1294
rect 41602 54 41736 82
rect 43810 82 43866 160
rect 43916 82 43944 1294
rect 44100 1222 44128 1906
rect 44560 1562 44588 1906
rect 44744 1834 44772 2314
rect 45020 2106 45048 2382
rect 45940 2106 45968 2382
rect 46670 2204 46978 2213
rect 46670 2202 46676 2204
rect 46732 2202 46756 2204
rect 46812 2202 46836 2204
rect 46892 2202 46916 2204
rect 46972 2202 46978 2204
rect 46732 2150 46734 2202
rect 46914 2150 46916 2202
rect 46670 2148 46676 2150
rect 46732 2148 46756 2150
rect 46812 2148 46836 2150
rect 46892 2148 46916 2150
rect 46972 2148 46978 2150
rect 46670 2139 46978 2148
rect 45008 2100 45060 2106
rect 45008 2042 45060 2048
rect 45928 2100 45980 2106
rect 45928 2042 45980 2048
rect 45652 1964 45704 1970
rect 45652 1906 45704 1912
rect 44732 1828 44784 1834
rect 44732 1770 44784 1776
rect 45664 1562 45692 1906
rect 44548 1556 44600 1562
rect 44548 1498 44600 1504
rect 45652 1556 45704 1562
rect 45652 1498 45704 1504
rect 46296 1352 46348 1358
rect 46296 1294 46348 1300
rect 44088 1216 44140 1222
rect 44088 1158 44140 1164
rect 43810 54 43944 82
rect 46018 82 46074 160
rect 46308 82 46336 1294
rect 46670 1116 46978 1125
rect 46670 1114 46676 1116
rect 46732 1114 46756 1116
rect 46812 1114 46836 1116
rect 46892 1114 46916 1116
rect 46972 1114 46978 1116
rect 46732 1062 46734 1114
rect 46914 1062 46916 1114
rect 46670 1060 46676 1062
rect 46732 1060 46756 1062
rect 46812 1060 46836 1062
rect 46892 1060 46916 1062
rect 46972 1060 46978 1062
rect 46670 1051 46978 1060
rect 46018 54 46336 82
rect 28354 0 28410 54
rect 30562 0 30618 54
rect 32770 0 32826 54
rect 34978 0 35034 54
rect 37186 0 37242 54
rect 39394 0 39450 54
rect 41602 0 41658 54
rect 43810 0 43866 54
rect 46018 0 46074 54
<< via2 >>
rect 2318 7792 2374 7848
rect 3238 6840 3294 6896
rect 6671 8186 6727 8188
rect 6751 8186 6807 8188
rect 6831 8186 6887 8188
rect 6911 8186 6967 8188
rect 6671 8134 6717 8186
rect 6717 8134 6727 8186
rect 6751 8134 6781 8186
rect 6781 8134 6793 8186
rect 6793 8134 6807 8186
rect 6831 8134 6845 8186
rect 6845 8134 6857 8186
rect 6857 8134 6887 8186
rect 6911 8134 6921 8186
rect 6921 8134 6967 8186
rect 6671 8132 6727 8134
rect 6751 8132 6807 8134
rect 6831 8132 6887 8134
rect 6911 8132 6967 8134
rect 6671 7098 6727 7100
rect 6751 7098 6807 7100
rect 6831 7098 6887 7100
rect 6911 7098 6967 7100
rect 6671 7046 6717 7098
rect 6717 7046 6727 7098
rect 6751 7046 6781 7098
rect 6781 7046 6793 7098
rect 6793 7046 6807 7098
rect 6831 7046 6845 7098
rect 6845 7046 6857 7098
rect 6857 7046 6887 7098
rect 6911 7046 6921 7098
rect 6921 7046 6967 7098
rect 6671 7044 6727 7046
rect 6751 7044 6807 7046
rect 6831 7044 6887 7046
rect 6911 7044 6967 7046
rect 12386 8730 12442 8732
rect 12466 8730 12522 8732
rect 12546 8730 12602 8732
rect 12626 8730 12682 8732
rect 12386 8678 12432 8730
rect 12432 8678 12442 8730
rect 12466 8678 12496 8730
rect 12496 8678 12508 8730
rect 12508 8678 12522 8730
rect 12546 8678 12560 8730
rect 12560 8678 12572 8730
rect 12572 8678 12602 8730
rect 12626 8678 12636 8730
rect 12636 8678 12682 8730
rect 12386 8676 12442 8678
rect 12466 8676 12522 8678
rect 12546 8676 12602 8678
rect 12626 8676 12682 8678
rect 11978 8200 12034 8256
rect 12990 9016 13046 9072
rect 13726 8880 13782 8936
rect 14646 9152 14702 9208
rect 14462 8356 14518 8392
rect 14462 8336 14464 8356
rect 14464 8336 14516 8356
rect 14516 8336 14518 8356
rect 14830 8508 14832 8528
rect 14832 8508 14884 8528
rect 14884 8508 14886 8528
rect 14830 8472 14886 8508
rect 12386 7642 12442 7644
rect 12466 7642 12522 7644
rect 12546 7642 12602 7644
rect 12626 7642 12682 7644
rect 12386 7590 12432 7642
rect 12432 7590 12442 7642
rect 12466 7590 12496 7642
rect 12496 7590 12508 7642
rect 12508 7590 12522 7642
rect 12546 7590 12560 7642
rect 12560 7590 12572 7642
rect 12572 7590 12602 7642
rect 12626 7590 12636 7642
rect 12636 7590 12682 7642
rect 12386 7588 12442 7590
rect 12466 7588 12522 7590
rect 12546 7588 12602 7590
rect 12626 7588 12682 7590
rect 14646 7520 14702 7576
rect 15106 7692 15108 7712
rect 15108 7692 15160 7712
rect 15160 7692 15162 7712
rect 15106 7656 15162 7692
rect 14830 7248 14886 7304
rect 16854 9560 16910 9616
rect 16210 8200 16266 8256
rect 17130 9424 17186 9480
rect 16946 7520 17002 7576
rect 16670 7384 16726 7440
rect 17866 9152 17922 9208
rect 17774 9016 17830 9072
rect 18101 8186 18157 8188
rect 18181 8186 18237 8188
rect 18261 8186 18317 8188
rect 18341 8186 18397 8188
rect 18101 8134 18147 8186
rect 18147 8134 18157 8186
rect 18181 8134 18211 8186
rect 18211 8134 18223 8186
rect 18223 8134 18237 8186
rect 18261 8134 18275 8186
rect 18275 8134 18287 8186
rect 18287 8134 18317 8186
rect 18341 8134 18351 8186
rect 18351 8134 18397 8186
rect 18101 8132 18157 8134
rect 18181 8132 18237 8134
rect 18261 8132 18317 8134
rect 18341 8132 18397 8134
rect 18510 8064 18566 8120
rect 17958 7928 18014 7984
rect 18970 9696 19026 9752
rect 19062 9560 19118 9616
rect 19798 9288 19854 9344
rect 19706 8608 19762 8664
rect 19338 8200 19394 8256
rect 19338 7692 19340 7712
rect 19340 7692 19392 7712
rect 19392 7692 19394 7712
rect 19338 7656 19394 7692
rect 18142 7520 18198 7576
rect 19982 9596 19984 9616
rect 19984 9596 20036 9616
rect 20036 9596 20038 9616
rect 19982 9560 20038 9596
rect 20074 9152 20130 9208
rect 20902 9560 20958 9616
rect 19982 7112 20038 7168
rect 18101 7098 18157 7100
rect 18181 7098 18237 7100
rect 18261 7098 18317 7100
rect 18341 7098 18397 7100
rect 18101 7046 18147 7098
rect 18147 7046 18157 7098
rect 18181 7046 18211 7098
rect 18211 7046 18223 7098
rect 18223 7046 18237 7098
rect 18261 7046 18275 7098
rect 18275 7046 18287 7098
rect 18287 7046 18317 7098
rect 18341 7046 18351 7098
rect 18351 7046 18397 7098
rect 18101 7044 18157 7046
rect 18181 7044 18237 7046
rect 18261 7044 18317 7046
rect 18341 7044 18397 7046
rect 12386 6554 12442 6556
rect 12466 6554 12522 6556
rect 12546 6554 12602 6556
rect 12626 6554 12682 6556
rect 12386 6502 12432 6554
rect 12432 6502 12442 6554
rect 12466 6502 12496 6554
rect 12496 6502 12508 6554
rect 12508 6502 12522 6554
rect 12546 6502 12560 6554
rect 12560 6502 12572 6554
rect 12572 6502 12602 6554
rect 12626 6502 12636 6554
rect 12636 6502 12682 6554
rect 12386 6500 12442 6502
rect 12466 6500 12522 6502
rect 12546 6500 12602 6502
rect 12626 6500 12682 6502
rect 21178 9424 21234 9480
rect 20902 8336 20958 8392
rect 21362 8744 21418 8800
rect 21638 9696 21694 9752
rect 21638 9036 21694 9072
rect 21638 9016 21640 9036
rect 21640 9016 21692 9036
rect 21692 9016 21694 9036
rect 21822 9288 21878 9344
rect 22282 9560 22338 9616
rect 21546 8336 21602 8392
rect 21362 8200 21418 8256
rect 22466 9052 22468 9072
rect 22468 9052 22520 9072
rect 22520 9052 22522 9072
rect 22466 9016 22522 9052
rect 21546 7520 21602 7576
rect 22650 9716 22706 9752
rect 22650 9696 22652 9716
rect 22652 9696 22704 9716
rect 22704 9696 22706 9716
rect 22742 8744 22798 8800
rect 22650 8628 22706 8664
rect 22650 8608 22652 8628
rect 22652 8608 22704 8628
rect 22704 8608 22706 8628
rect 24030 9288 24086 9344
rect 23816 8730 23872 8732
rect 23896 8730 23952 8732
rect 23976 8730 24032 8732
rect 24056 8730 24112 8732
rect 23816 8678 23862 8730
rect 23862 8678 23872 8730
rect 23896 8678 23926 8730
rect 23926 8678 23938 8730
rect 23938 8678 23952 8730
rect 23976 8678 23990 8730
rect 23990 8678 24002 8730
rect 24002 8678 24032 8730
rect 24056 8678 24066 8730
rect 24066 8678 24112 8730
rect 23816 8676 23872 8678
rect 23896 8676 23952 8678
rect 23976 8676 24032 8678
rect 24056 8676 24112 8678
rect 22834 7656 22890 7712
rect 23386 7384 23442 7440
rect 23754 8372 23756 8392
rect 23756 8372 23808 8392
rect 23808 8372 23810 8392
rect 23754 8336 23810 8372
rect 23846 8200 23902 8256
rect 24766 9460 24768 9480
rect 24768 9460 24820 9480
rect 24820 9460 24822 9480
rect 24766 9424 24822 9460
rect 24674 9152 24730 9208
rect 24398 8336 24454 8392
rect 23816 7642 23872 7644
rect 23896 7642 23952 7644
rect 23976 7642 24032 7644
rect 24056 7642 24112 7644
rect 23816 7590 23862 7642
rect 23862 7590 23872 7642
rect 23896 7590 23926 7642
rect 23926 7590 23938 7642
rect 23938 7590 23952 7642
rect 23976 7590 23990 7642
rect 23990 7590 24002 7642
rect 24002 7590 24032 7642
rect 24056 7590 24066 7642
rect 24066 7590 24112 7642
rect 23816 7588 23872 7590
rect 23896 7588 23952 7590
rect 23976 7588 24032 7590
rect 24056 7588 24112 7590
rect 23816 6554 23872 6556
rect 23896 6554 23952 6556
rect 23976 6554 24032 6556
rect 24056 6554 24112 6556
rect 23816 6502 23862 6554
rect 23862 6502 23872 6554
rect 23896 6502 23926 6554
rect 23926 6502 23938 6554
rect 23938 6502 23952 6554
rect 23976 6502 23990 6554
rect 23990 6502 24002 6554
rect 24002 6502 24032 6554
rect 24056 6502 24066 6554
rect 24066 6502 24112 6554
rect 23816 6500 23872 6502
rect 23896 6500 23952 6502
rect 23976 6500 24032 6502
rect 24056 6500 24112 6502
rect 25410 8472 25466 8528
rect 27710 9560 27766 9616
rect 26790 7692 26792 7712
rect 26792 7692 26844 7712
rect 26844 7692 26846 7712
rect 26790 7656 26846 7692
rect 28078 8880 28134 8936
rect 28354 9696 28410 9752
rect 28170 8336 28226 8392
rect 28262 8200 28318 8256
rect 27986 7112 28042 7168
rect 29531 8186 29587 8188
rect 29611 8186 29667 8188
rect 29691 8186 29747 8188
rect 29771 8186 29827 8188
rect 29531 8134 29577 8186
rect 29577 8134 29587 8186
rect 29611 8134 29641 8186
rect 29641 8134 29653 8186
rect 29653 8134 29667 8186
rect 29691 8134 29705 8186
rect 29705 8134 29717 8186
rect 29717 8134 29747 8186
rect 29771 8134 29781 8186
rect 29781 8134 29827 8186
rect 29531 8132 29587 8134
rect 29611 8132 29667 8134
rect 29691 8132 29747 8134
rect 29771 8132 29827 8134
rect 29182 7248 29238 7304
rect 29531 7098 29587 7100
rect 29611 7098 29667 7100
rect 29691 7098 29747 7100
rect 29771 7098 29827 7100
rect 29531 7046 29577 7098
rect 29577 7046 29587 7098
rect 29611 7046 29641 7098
rect 29641 7046 29653 7098
rect 29653 7046 29667 7098
rect 29691 7046 29705 7098
rect 29705 7046 29717 7098
rect 29717 7046 29747 7098
rect 29771 7046 29781 7098
rect 29781 7046 29827 7098
rect 29531 7044 29587 7046
rect 29611 7044 29667 7046
rect 29691 7044 29747 7046
rect 29771 7044 29827 7046
rect 26238 6840 26294 6896
rect 6671 6010 6727 6012
rect 6751 6010 6807 6012
rect 6831 6010 6887 6012
rect 6911 6010 6967 6012
rect 6671 5958 6717 6010
rect 6717 5958 6727 6010
rect 6751 5958 6781 6010
rect 6781 5958 6793 6010
rect 6793 5958 6807 6010
rect 6831 5958 6845 6010
rect 6845 5958 6857 6010
rect 6857 5958 6887 6010
rect 6911 5958 6921 6010
rect 6921 5958 6967 6010
rect 6671 5956 6727 5958
rect 6751 5956 6807 5958
rect 6831 5956 6887 5958
rect 6911 5956 6967 5958
rect 18101 6010 18157 6012
rect 18181 6010 18237 6012
rect 18261 6010 18317 6012
rect 18341 6010 18397 6012
rect 18101 5958 18147 6010
rect 18147 5958 18157 6010
rect 18181 5958 18211 6010
rect 18211 5958 18223 6010
rect 18223 5958 18237 6010
rect 18261 5958 18275 6010
rect 18275 5958 18287 6010
rect 18287 5958 18317 6010
rect 18341 5958 18351 6010
rect 18351 5958 18397 6010
rect 18101 5956 18157 5958
rect 18181 5956 18237 5958
rect 18261 5956 18317 5958
rect 18341 5956 18397 5958
rect 12386 5466 12442 5468
rect 12466 5466 12522 5468
rect 12546 5466 12602 5468
rect 12626 5466 12682 5468
rect 12386 5414 12432 5466
rect 12432 5414 12442 5466
rect 12466 5414 12496 5466
rect 12496 5414 12508 5466
rect 12508 5414 12522 5466
rect 12546 5414 12560 5466
rect 12560 5414 12572 5466
rect 12572 5414 12602 5466
rect 12626 5414 12636 5466
rect 12636 5414 12682 5466
rect 12386 5412 12442 5414
rect 12466 5412 12522 5414
rect 12546 5412 12602 5414
rect 12626 5412 12682 5414
rect 23816 5466 23872 5468
rect 23896 5466 23952 5468
rect 23976 5466 24032 5468
rect 24056 5466 24112 5468
rect 23816 5414 23862 5466
rect 23862 5414 23872 5466
rect 23896 5414 23926 5466
rect 23926 5414 23938 5466
rect 23938 5414 23952 5466
rect 23976 5414 23990 5466
rect 23990 5414 24002 5466
rect 24002 5414 24032 5466
rect 24056 5414 24066 5466
rect 24066 5414 24112 5466
rect 23816 5412 23872 5414
rect 23896 5412 23952 5414
rect 23976 5412 24032 5414
rect 24056 5412 24112 5414
rect 6671 4922 6727 4924
rect 6751 4922 6807 4924
rect 6831 4922 6887 4924
rect 6911 4922 6967 4924
rect 6671 4870 6717 4922
rect 6717 4870 6727 4922
rect 6751 4870 6781 4922
rect 6781 4870 6793 4922
rect 6793 4870 6807 4922
rect 6831 4870 6845 4922
rect 6845 4870 6857 4922
rect 6857 4870 6887 4922
rect 6911 4870 6921 4922
rect 6921 4870 6967 4922
rect 6671 4868 6727 4870
rect 6751 4868 6807 4870
rect 6831 4868 6887 4870
rect 6911 4868 6967 4870
rect 18101 4922 18157 4924
rect 18181 4922 18237 4924
rect 18261 4922 18317 4924
rect 18341 4922 18397 4924
rect 18101 4870 18147 4922
rect 18147 4870 18157 4922
rect 18181 4870 18211 4922
rect 18211 4870 18223 4922
rect 18223 4870 18237 4922
rect 18261 4870 18275 4922
rect 18275 4870 18287 4922
rect 18287 4870 18317 4922
rect 18341 4870 18351 4922
rect 18351 4870 18397 4922
rect 18101 4868 18157 4870
rect 18181 4868 18237 4870
rect 18261 4868 18317 4870
rect 18341 4868 18397 4870
rect 12386 4378 12442 4380
rect 12466 4378 12522 4380
rect 12546 4378 12602 4380
rect 12626 4378 12682 4380
rect 12386 4326 12432 4378
rect 12432 4326 12442 4378
rect 12466 4326 12496 4378
rect 12496 4326 12508 4378
rect 12508 4326 12522 4378
rect 12546 4326 12560 4378
rect 12560 4326 12572 4378
rect 12572 4326 12602 4378
rect 12626 4326 12636 4378
rect 12636 4326 12682 4378
rect 12386 4324 12442 4326
rect 12466 4324 12522 4326
rect 12546 4324 12602 4326
rect 12626 4324 12682 4326
rect 23816 4378 23872 4380
rect 23896 4378 23952 4380
rect 23976 4378 24032 4380
rect 24056 4378 24112 4380
rect 23816 4326 23862 4378
rect 23862 4326 23872 4378
rect 23896 4326 23926 4378
rect 23926 4326 23938 4378
rect 23938 4326 23952 4378
rect 23976 4326 23990 4378
rect 23990 4326 24002 4378
rect 24002 4326 24032 4378
rect 24056 4326 24066 4378
rect 24066 4326 24112 4378
rect 23816 4324 23872 4326
rect 23896 4324 23952 4326
rect 23976 4324 24032 4326
rect 24056 4324 24112 4326
rect 6671 3834 6727 3836
rect 6751 3834 6807 3836
rect 6831 3834 6887 3836
rect 6911 3834 6967 3836
rect 6671 3782 6717 3834
rect 6717 3782 6727 3834
rect 6751 3782 6781 3834
rect 6781 3782 6793 3834
rect 6793 3782 6807 3834
rect 6831 3782 6845 3834
rect 6845 3782 6857 3834
rect 6857 3782 6887 3834
rect 6911 3782 6921 3834
rect 6921 3782 6967 3834
rect 6671 3780 6727 3782
rect 6751 3780 6807 3782
rect 6831 3780 6887 3782
rect 6911 3780 6967 3782
rect 18101 3834 18157 3836
rect 18181 3834 18237 3836
rect 18261 3834 18317 3836
rect 18341 3834 18397 3836
rect 18101 3782 18147 3834
rect 18147 3782 18157 3834
rect 18181 3782 18211 3834
rect 18211 3782 18223 3834
rect 18223 3782 18237 3834
rect 18261 3782 18275 3834
rect 18275 3782 18287 3834
rect 18287 3782 18317 3834
rect 18341 3782 18351 3834
rect 18351 3782 18397 3834
rect 18101 3780 18157 3782
rect 18181 3780 18237 3782
rect 18261 3780 18317 3782
rect 18341 3780 18397 3782
rect 12386 3290 12442 3292
rect 12466 3290 12522 3292
rect 12546 3290 12602 3292
rect 12626 3290 12682 3292
rect 12386 3238 12432 3290
rect 12432 3238 12442 3290
rect 12466 3238 12496 3290
rect 12496 3238 12508 3290
rect 12508 3238 12522 3290
rect 12546 3238 12560 3290
rect 12560 3238 12572 3290
rect 12572 3238 12602 3290
rect 12626 3238 12636 3290
rect 12636 3238 12682 3290
rect 12386 3236 12442 3238
rect 12466 3236 12522 3238
rect 12546 3236 12602 3238
rect 12626 3236 12682 3238
rect 6671 2746 6727 2748
rect 6751 2746 6807 2748
rect 6831 2746 6887 2748
rect 6911 2746 6967 2748
rect 6671 2694 6717 2746
rect 6717 2694 6727 2746
rect 6751 2694 6781 2746
rect 6781 2694 6793 2746
rect 6793 2694 6807 2746
rect 6831 2694 6845 2746
rect 6845 2694 6857 2746
rect 6857 2694 6887 2746
rect 6911 2694 6921 2746
rect 6921 2694 6967 2746
rect 6671 2692 6727 2694
rect 6751 2692 6807 2694
rect 6831 2692 6887 2694
rect 6911 2692 6967 2694
rect 18101 2746 18157 2748
rect 18181 2746 18237 2748
rect 18261 2746 18317 2748
rect 18341 2746 18397 2748
rect 18101 2694 18147 2746
rect 18147 2694 18157 2746
rect 18181 2694 18211 2746
rect 18211 2694 18223 2746
rect 18223 2694 18237 2746
rect 18261 2694 18275 2746
rect 18275 2694 18287 2746
rect 18287 2694 18317 2746
rect 18341 2694 18351 2746
rect 18351 2694 18397 2746
rect 18101 2692 18157 2694
rect 18181 2692 18237 2694
rect 18261 2692 18317 2694
rect 18341 2692 18397 2694
rect 23816 3290 23872 3292
rect 23896 3290 23952 3292
rect 23976 3290 24032 3292
rect 24056 3290 24112 3292
rect 23816 3238 23862 3290
rect 23862 3238 23872 3290
rect 23896 3238 23926 3290
rect 23926 3238 23938 3290
rect 23938 3238 23952 3290
rect 23976 3238 23990 3290
rect 23990 3238 24002 3290
rect 24002 3238 24032 3290
rect 24056 3238 24066 3290
rect 24066 3238 24112 3290
rect 23816 3236 23872 3238
rect 23896 3236 23952 3238
rect 23976 3236 24032 3238
rect 24056 3236 24112 3238
rect 12386 2202 12442 2204
rect 12466 2202 12522 2204
rect 12546 2202 12602 2204
rect 12626 2202 12682 2204
rect 12386 2150 12432 2202
rect 12432 2150 12442 2202
rect 12466 2150 12496 2202
rect 12496 2150 12508 2202
rect 12508 2150 12522 2202
rect 12546 2150 12560 2202
rect 12560 2150 12572 2202
rect 12572 2150 12602 2202
rect 12626 2150 12636 2202
rect 12636 2150 12682 2202
rect 12386 2148 12442 2150
rect 12466 2148 12522 2150
rect 12546 2148 12602 2150
rect 12626 2148 12682 2150
rect 6671 1658 6727 1660
rect 6751 1658 6807 1660
rect 6831 1658 6887 1660
rect 6911 1658 6967 1660
rect 6671 1606 6717 1658
rect 6717 1606 6727 1658
rect 6751 1606 6781 1658
rect 6781 1606 6793 1658
rect 6793 1606 6807 1658
rect 6831 1606 6845 1658
rect 6845 1606 6857 1658
rect 6857 1606 6887 1658
rect 6911 1606 6921 1658
rect 6921 1606 6967 1658
rect 6671 1604 6727 1606
rect 6751 1604 6807 1606
rect 6831 1604 6887 1606
rect 6911 1604 6967 1606
rect 18101 1658 18157 1660
rect 18181 1658 18237 1660
rect 18261 1658 18317 1660
rect 18341 1658 18397 1660
rect 18101 1606 18147 1658
rect 18147 1606 18157 1658
rect 18181 1606 18211 1658
rect 18211 1606 18223 1658
rect 18223 1606 18237 1658
rect 18261 1606 18275 1658
rect 18275 1606 18287 1658
rect 18287 1606 18317 1658
rect 18341 1606 18351 1658
rect 18351 1606 18397 1658
rect 18101 1604 18157 1606
rect 18181 1604 18237 1606
rect 18261 1604 18317 1606
rect 18341 1604 18397 1606
rect 12386 1114 12442 1116
rect 12466 1114 12522 1116
rect 12546 1114 12602 1116
rect 12626 1114 12682 1116
rect 12386 1062 12432 1114
rect 12432 1062 12442 1114
rect 12466 1062 12496 1114
rect 12496 1062 12508 1114
rect 12508 1062 12522 1114
rect 12546 1062 12560 1114
rect 12560 1062 12572 1114
rect 12572 1062 12602 1114
rect 12626 1062 12636 1114
rect 12636 1062 12682 1114
rect 12386 1060 12442 1062
rect 12466 1060 12522 1062
rect 12546 1060 12602 1062
rect 12626 1060 12682 1062
rect 23816 2202 23872 2204
rect 23896 2202 23952 2204
rect 23976 2202 24032 2204
rect 24056 2202 24112 2204
rect 23816 2150 23862 2202
rect 23862 2150 23872 2202
rect 23896 2150 23926 2202
rect 23926 2150 23938 2202
rect 23938 2150 23952 2202
rect 23976 2150 23990 2202
rect 23990 2150 24002 2202
rect 24002 2150 24032 2202
rect 24056 2150 24066 2202
rect 24066 2150 24112 2202
rect 23816 2148 23872 2150
rect 23896 2148 23952 2150
rect 23976 2148 24032 2150
rect 24056 2148 24112 2150
rect 29531 6010 29587 6012
rect 29611 6010 29667 6012
rect 29691 6010 29747 6012
rect 29771 6010 29827 6012
rect 29531 5958 29577 6010
rect 29577 5958 29587 6010
rect 29611 5958 29641 6010
rect 29641 5958 29653 6010
rect 29653 5958 29667 6010
rect 29691 5958 29705 6010
rect 29705 5958 29717 6010
rect 29717 5958 29747 6010
rect 29771 5958 29781 6010
rect 29781 5958 29827 6010
rect 29531 5956 29587 5958
rect 29611 5956 29667 5958
rect 29691 5956 29747 5958
rect 29771 5956 29827 5958
rect 29531 4922 29587 4924
rect 29611 4922 29667 4924
rect 29691 4922 29747 4924
rect 29771 4922 29827 4924
rect 29531 4870 29577 4922
rect 29577 4870 29587 4922
rect 29611 4870 29641 4922
rect 29641 4870 29653 4922
rect 29653 4870 29667 4922
rect 29691 4870 29705 4922
rect 29705 4870 29717 4922
rect 29717 4870 29747 4922
rect 29771 4870 29781 4922
rect 29781 4870 29827 4922
rect 29531 4868 29587 4870
rect 29611 4868 29667 4870
rect 29691 4868 29747 4870
rect 29771 4868 29827 4870
rect 23816 1114 23872 1116
rect 23896 1114 23952 1116
rect 23976 1114 24032 1116
rect 24056 1114 24112 1116
rect 23816 1062 23862 1114
rect 23862 1062 23872 1114
rect 23896 1062 23926 1114
rect 23926 1062 23938 1114
rect 23938 1062 23952 1114
rect 23976 1062 23990 1114
rect 23990 1062 24002 1114
rect 24002 1062 24032 1114
rect 24056 1062 24066 1114
rect 24066 1062 24112 1114
rect 23816 1060 23872 1062
rect 23896 1060 23952 1062
rect 23976 1060 24032 1062
rect 24056 1060 24112 1062
rect 29531 3834 29587 3836
rect 29611 3834 29667 3836
rect 29691 3834 29747 3836
rect 29771 3834 29827 3836
rect 29531 3782 29577 3834
rect 29577 3782 29587 3834
rect 29611 3782 29641 3834
rect 29641 3782 29653 3834
rect 29653 3782 29667 3834
rect 29691 3782 29705 3834
rect 29705 3782 29717 3834
rect 29717 3782 29747 3834
rect 29771 3782 29781 3834
rect 29781 3782 29827 3834
rect 29531 3780 29587 3782
rect 29611 3780 29667 3782
rect 29691 3780 29747 3782
rect 29771 3780 29827 3782
rect 29531 2746 29587 2748
rect 29611 2746 29667 2748
rect 29691 2746 29747 2748
rect 29771 2746 29827 2748
rect 29531 2694 29577 2746
rect 29577 2694 29587 2746
rect 29611 2694 29641 2746
rect 29641 2694 29653 2746
rect 29653 2694 29667 2746
rect 29691 2694 29705 2746
rect 29705 2694 29717 2746
rect 29717 2694 29747 2746
rect 29771 2694 29781 2746
rect 29781 2694 29827 2746
rect 29531 2692 29587 2694
rect 29611 2692 29667 2694
rect 29691 2692 29747 2694
rect 29771 2692 29827 2694
rect 35246 8730 35302 8732
rect 35326 8730 35382 8732
rect 35406 8730 35462 8732
rect 35486 8730 35542 8732
rect 35246 8678 35292 8730
rect 35292 8678 35302 8730
rect 35326 8678 35356 8730
rect 35356 8678 35368 8730
rect 35368 8678 35382 8730
rect 35406 8678 35420 8730
rect 35420 8678 35432 8730
rect 35432 8678 35462 8730
rect 35486 8678 35496 8730
rect 35496 8678 35542 8730
rect 35246 8676 35302 8678
rect 35326 8676 35382 8678
rect 35406 8676 35462 8678
rect 35486 8676 35542 8678
rect 35070 8064 35126 8120
rect 35806 7928 35862 7984
rect 35246 7642 35302 7644
rect 35326 7642 35382 7644
rect 35406 7642 35462 7644
rect 35486 7642 35542 7644
rect 35246 7590 35292 7642
rect 35292 7590 35302 7642
rect 35326 7590 35356 7642
rect 35356 7590 35368 7642
rect 35368 7590 35382 7642
rect 35406 7590 35420 7642
rect 35420 7590 35432 7642
rect 35432 7590 35462 7642
rect 35486 7590 35496 7642
rect 35496 7590 35542 7642
rect 35246 7588 35302 7590
rect 35326 7588 35382 7590
rect 35406 7588 35462 7590
rect 35486 7588 35542 7590
rect 35246 6554 35302 6556
rect 35326 6554 35382 6556
rect 35406 6554 35462 6556
rect 35486 6554 35542 6556
rect 35246 6502 35292 6554
rect 35292 6502 35302 6554
rect 35326 6502 35356 6554
rect 35356 6502 35368 6554
rect 35368 6502 35382 6554
rect 35406 6502 35420 6554
rect 35420 6502 35432 6554
rect 35432 6502 35462 6554
rect 35486 6502 35496 6554
rect 35496 6502 35542 6554
rect 35246 6500 35302 6502
rect 35326 6500 35382 6502
rect 35406 6500 35462 6502
rect 35486 6500 35542 6502
rect 35246 5466 35302 5468
rect 35326 5466 35382 5468
rect 35406 5466 35462 5468
rect 35486 5466 35542 5468
rect 35246 5414 35292 5466
rect 35292 5414 35302 5466
rect 35326 5414 35356 5466
rect 35356 5414 35368 5466
rect 35368 5414 35382 5466
rect 35406 5414 35420 5466
rect 35420 5414 35432 5466
rect 35432 5414 35462 5466
rect 35486 5414 35496 5466
rect 35496 5414 35542 5466
rect 35246 5412 35302 5414
rect 35326 5412 35382 5414
rect 35406 5412 35462 5414
rect 35486 5412 35542 5414
rect 35246 4378 35302 4380
rect 35326 4378 35382 4380
rect 35406 4378 35462 4380
rect 35486 4378 35542 4380
rect 35246 4326 35292 4378
rect 35292 4326 35302 4378
rect 35326 4326 35356 4378
rect 35356 4326 35368 4378
rect 35368 4326 35382 4378
rect 35406 4326 35420 4378
rect 35420 4326 35432 4378
rect 35432 4326 35462 4378
rect 35486 4326 35496 4378
rect 35496 4326 35542 4378
rect 35246 4324 35302 4326
rect 35326 4324 35382 4326
rect 35406 4324 35462 4326
rect 35486 4324 35542 4326
rect 35246 3290 35302 3292
rect 35326 3290 35382 3292
rect 35406 3290 35462 3292
rect 35486 3290 35542 3292
rect 35246 3238 35292 3290
rect 35292 3238 35302 3290
rect 35326 3238 35356 3290
rect 35356 3238 35368 3290
rect 35368 3238 35382 3290
rect 35406 3238 35420 3290
rect 35420 3238 35432 3290
rect 35432 3238 35462 3290
rect 35486 3238 35496 3290
rect 35496 3238 35542 3290
rect 35246 3236 35302 3238
rect 35326 3236 35382 3238
rect 35406 3236 35462 3238
rect 35486 3236 35542 3238
rect 35246 2202 35302 2204
rect 35326 2202 35382 2204
rect 35406 2202 35462 2204
rect 35486 2202 35542 2204
rect 35246 2150 35292 2202
rect 35292 2150 35302 2202
rect 35326 2150 35356 2202
rect 35356 2150 35368 2202
rect 35368 2150 35382 2202
rect 35406 2150 35420 2202
rect 35420 2150 35432 2202
rect 35432 2150 35462 2202
rect 35486 2150 35496 2202
rect 35496 2150 35542 2202
rect 35246 2148 35302 2150
rect 35326 2148 35382 2150
rect 35406 2148 35462 2150
rect 35486 2148 35542 2150
rect 29531 1658 29587 1660
rect 29611 1658 29667 1660
rect 29691 1658 29747 1660
rect 29771 1658 29827 1660
rect 29531 1606 29577 1658
rect 29577 1606 29587 1658
rect 29611 1606 29641 1658
rect 29641 1606 29653 1658
rect 29653 1606 29667 1658
rect 29691 1606 29705 1658
rect 29705 1606 29717 1658
rect 29717 1606 29747 1658
rect 29771 1606 29781 1658
rect 29781 1606 29827 1658
rect 29531 1604 29587 1606
rect 29611 1604 29667 1606
rect 29691 1604 29747 1606
rect 29771 1604 29827 1606
rect 38750 7384 38806 7440
rect 40961 8186 41017 8188
rect 41041 8186 41097 8188
rect 41121 8186 41177 8188
rect 41201 8186 41257 8188
rect 40961 8134 41007 8186
rect 41007 8134 41017 8186
rect 41041 8134 41071 8186
rect 41071 8134 41083 8186
rect 41083 8134 41097 8186
rect 41121 8134 41135 8186
rect 41135 8134 41147 8186
rect 41147 8134 41177 8186
rect 41201 8134 41211 8186
rect 41211 8134 41257 8186
rect 40961 8132 41017 8134
rect 41041 8132 41097 8134
rect 41121 8132 41177 8134
rect 41201 8132 41257 8134
rect 40961 7098 41017 7100
rect 41041 7098 41097 7100
rect 41121 7098 41177 7100
rect 41201 7098 41257 7100
rect 40961 7046 41007 7098
rect 41007 7046 41017 7098
rect 41041 7046 41071 7098
rect 41071 7046 41083 7098
rect 41083 7046 41097 7098
rect 41121 7046 41135 7098
rect 41135 7046 41147 7098
rect 41147 7046 41177 7098
rect 41201 7046 41211 7098
rect 41211 7046 41257 7098
rect 40961 7044 41017 7046
rect 41041 7044 41097 7046
rect 41121 7044 41177 7046
rect 41201 7044 41257 7046
rect 40961 6010 41017 6012
rect 41041 6010 41097 6012
rect 41121 6010 41177 6012
rect 41201 6010 41257 6012
rect 40961 5958 41007 6010
rect 41007 5958 41017 6010
rect 41041 5958 41071 6010
rect 41071 5958 41083 6010
rect 41083 5958 41097 6010
rect 41121 5958 41135 6010
rect 41135 5958 41147 6010
rect 41147 5958 41177 6010
rect 41201 5958 41211 6010
rect 41211 5958 41257 6010
rect 40961 5956 41017 5958
rect 41041 5956 41097 5958
rect 41121 5956 41177 5958
rect 41201 5956 41257 5958
rect 40961 4922 41017 4924
rect 41041 4922 41097 4924
rect 41121 4922 41177 4924
rect 41201 4922 41257 4924
rect 40961 4870 41007 4922
rect 41007 4870 41017 4922
rect 41041 4870 41071 4922
rect 41071 4870 41083 4922
rect 41083 4870 41097 4922
rect 41121 4870 41135 4922
rect 41135 4870 41147 4922
rect 41147 4870 41177 4922
rect 41201 4870 41211 4922
rect 41211 4870 41257 4922
rect 40961 4868 41017 4870
rect 41041 4868 41097 4870
rect 41121 4868 41177 4870
rect 41201 4868 41257 4870
rect 40961 3834 41017 3836
rect 41041 3834 41097 3836
rect 41121 3834 41177 3836
rect 41201 3834 41257 3836
rect 40961 3782 41007 3834
rect 41007 3782 41017 3834
rect 41041 3782 41071 3834
rect 41071 3782 41083 3834
rect 41083 3782 41097 3834
rect 41121 3782 41135 3834
rect 41135 3782 41147 3834
rect 41147 3782 41177 3834
rect 41201 3782 41211 3834
rect 41211 3782 41257 3834
rect 40961 3780 41017 3782
rect 41041 3780 41097 3782
rect 41121 3780 41177 3782
rect 41201 3780 41257 3782
rect 40961 2746 41017 2748
rect 41041 2746 41097 2748
rect 41121 2746 41177 2748
rect 41201 2746 41257 2748
rect 40961 2694 41007 2746
rect 41007 2694 41017 2746
rect 41041 2694 41071 2746
rect 41071 2694 41083 2746
rect 41083 2694 41097 2746
rect 41121 2694 41135 2746
rect 41135 2694 41147 2746
rect 41147 2694 41177 2746
rect 41201 2694 41211 2746
rect 41211 2694 41257 2746
rect 40961 2692 41017 2694
rect 41041 2692 41097 2694
rect 41121 2692 41177 2694
rect 41201 2692 41257 2694
rect 46676 8730 46732 8732
rect 46756 8730 46812 8732
rect 46836 8730 46892 8732
rect 46916 8730 46972 8732
rect 46676 8678 46722 8730
rect 46722 8678 46732 8730
rect 46756 8678 46786 8730
rect 46786 8678 46798 8730
rect 46798 8678 46812 8730
rect 46836 8678 46850 8730
rect 46850 8678 46862 8730
rect 46862 8678 46892 8730
rect 46916 8678 46926 8730
rect 46926 8678 46972 8730
rect 46676 8676 46732 8678
rect 46756 8676 46812 8678
rect 46836 8676 46892 8678
rect 46916 8676 46972 8678
rect 46676 7642 46732 7644
rect 46756 7642 46812 7644
rect 46836 7642 46892 7644
rect 46916 7642 46972 7644
rect 46676 7590 46722 7642
rect 46722 7590 46732 7642
rect 46756 7590 46786 7642
rect 46786 7590 46798 7642
rect 46798 7590 46812 7642
rect 46836 7590 46850 7642
rect 46850 7590 46862 7642
rect 46862 7590 46892 7642
rect 46916 7590 46926 7642
rect 46926 7590 46972 7642
rect 46676 7588 46732 7590
rect 46756 7588 46812 7590
rect 46836 7588 46892 7590
rect 46916 7588 46972 7590
rect 46676 6554 46732 6556
rect 46756 6554 46812 6556
rect 46836 6554 46892 6556
rect 46916 6554 46972 6556
rect 46676 6502 46722 6554
rect 46722 6502 46732 6554
rect 46756 6502 46786 6554
rect 46786 6502 46798 6554
rect 46798 6502 46812 6554
rect 46836 6502 46850 6554
rect 46850 6502 46862 6554
rect 46862 6502 46892 6554
rect 46916 6502 46926 6554
rect 46926 6502 46972 6554
rect 46676 6500 46732 6502
rect 46756 6500 46812 6502
rect 46836 6500 46892 6502
rect 46916 6500 46972 6502
rect 46676 5466 46732 5468
rect 46756 5466 46812 5468
rect 46836 5466 46892 5468
rect 46916 5466 46972 5468
rect 46676 5414 46722 5466
rect 46722 5414 46732 5466
rect 46756 5414 46786 5466
rect 46786 5414 46798 5466
rect 46798 5414 46812 5466
rect 46836 5414 46850 5466
rect 46850 5414 46862 5466
rect 46862 5414 46892 5466
rect 46916 5414 46926 5466
rect 46926 5414 46972 5466
rect 46676 5412 46732 5414
rect 46756 5412 46812 5414
rect 46836 5412 46892 5414
rect 46916 5412 46972 5414
rect 46676 4378 46732 4380
rect 46756 4378 46812 4380
rect 46836 4378 46892 4380
rect 46916 4378 46972 4380
rect 46676 4326 46722 4378
rect 46722 4326 46732 4378
rect 46756 4326 46786 4378
rect 46786 4326 46798 4378
rect 46798 4326 46812 4378
rect 46836 4326 46850 4378
rect 46850 4326 46862 4378
rect 46862 4326 46892 4378
rect 46916 4326 46926 4378
rect 46926 4326 46972 4378
rect 46676 4324 46732 4326
rect 46756 4324 46812 4326
rect 46836 4324 46892 4326
rect 46916 4324 46972 4326
rect 46676 3290 46732 3292
rect 46756 3290 46812 3292
rect 46836 3290 46892 3292
rect 46916 3290 46972 3292
rect 46676 3238 46722 3290
rect 46722 3238 46732 3290
rect 46756 3238 46786 3290
rect 46786 3238 46798 3290
rect 46798 3238 46812 3290
rect 46836 3238 46850 3290
rect 46850 3238 46862 3290
rect 46862 3238 46892 3290
rect 46916 3238 46926 3290
rect 46926 3238 46972 3290
rect 46676 3236 46732 3238
rect 46756 3236 46812 3238
rect 46836 3236 46892 3238
rect 46916 3236 46972 3238
rect 40961 1658 41017 1660
rect 41041 1658 41097 1660
rect 41121 1658 41177 1660
rect 41201 1658 41257 1660
rect 40961 1606 41007 1658
rect 41007 1606 41017 1658
rect 41041 1606 41071 1658
rect 41071 1606 41083 1658
rect 41083 1606 41097 1658
rect 41121 1606 41135 1658
rect 41135 1606 41147 1658
rect 41147 1606 41177 1658
rect 41201 1606 41211 1658
rect 41211 1606 41257 1658
rect 40961 1604 41017 1606
rect 41041 1604 41097 1606
rect 41121 1604 41177 1606
rect 41201 1604 41257 1606
rect 35246 1114 35302 1116
rect 35326 1114 35382 1116
rect 35406 1114 35462 1116
rect 35486 1114 35542 1116
rect 35246 1062 35292 1114
rect 35292 1062 35302 1114
rect 35326 1062 35356 1114
rect 35356 1062 35368 1114
rect 35368 1062 35382 1114
rect 35406 1062 35420 1114
rect 35420 1062 35432 1114
rect 35432 1062 35462 1114
rect 35486 1062 35496 1114
rect 35496 1062 35542 1114
rect 35246 1060 35302 1062
rect 35326 1060 35382 1062
rect 35406 1060 35462 1062
rect 35486 1060 35542 1062
rect 46676 2202 46732 2204
rect 46756 2202 46812 2204
rect 46836 2202 46892 2204
rect 46916 2202 46972 2204
rect 46676 2150 46722 2202
rect 46722 2150 46732 2202
rect 46756 2150 46786 2202
rect 46786 2150 46798 2202
rect 46798 2150 46812 2202
rect 46836 2150 46850 2202
rect 46850 2150 46862 2202
rect 46862 2150 46892 2202
rect 46916 2150 46926 2202
rect 46926 2150 46972 2202
rect 46676 2148 46732 2150
rect 46756 2148 46812 2150
rect 46836 2148 46892 2150
rect 46916 2148 46972 2150
rect 46676 1114 46732 1116
rect 46756 1114 46812 1116
rect 46836 1114 46892 1116
rect 46916 1114 46972 1116
rect 46676 1062 46722 1114
rect 46722 1062 46732 1114
rect 46756 1062 46786 1114
rect 46786 1062 46798 1114
rect 46798 1062 46812 1114
rect 46836 1062 46850 1114
rect 46850 1062 46862 1114
rect 46862 1062 46892 1114
rect 46916 1062 46926 1114
rect 46926 1062 46972 1114
rect 46676 1060 46732 1062
rect 46756 1060 46812 1062
rect 46836 1060 46892 1062
rect 46916 1060 46972 1062
<< metal3 >>
rect 19290 9830 22892 9890
rect 18965 9754 19031 9757
rect 19290 9754 19350 9830
rect 18965 9752 19350 9754
rect 18965 9696 18970 9752
rect 19026 9696 19350 9752
rect 18965 9694 19350 9696
rect 21633 9754 21699 9757
rect 22645 9754 22711 9757
rect 21633 9752 22711 9754
rect 21633 9696 21638 9752
rect 21694 9696 22650 9752
rect 22706 9696 22711 9752
rect 21633 9694 22711 9696
rect 22832 9754 22892 9830
rect 28349 9754 28415 9757
rect 22832 9752 28415 9754
rect 22832 9696 28354 9752
rect 28410 9696 28415 9752
rect 22832 9694 28415 9696
rect 18965 9691 19031 9694
rect 21633 9691 21699 9694
rect 22645 9691 22711 9694
rect 28349 9691 28415 9694
rect 16849 9618 16915 9621
rect 19057 9618 19123 9621
rect 16849 9616 19123 9618
rect 16849 9560 16854 9616
rect 16910 9560 19062 9616
rect 19118 9560 19123 9616
rect 16849 9558 19123 9560
rect 16849 9555 16915 9558
rect 19057 9555 19123 9558
rect 19977 9618 20043 9621
rect 20897 9618 20963 9621
rect 19977 9616 20963 9618
rect 19977 9560 19982 9616
rect 20038 9560 20902 9616
rect 20958 9560 20963 9616
rect 19977 9558 20963 9560
rect 19977 9555 20043 9558
rect 20897 9555 20963 9558
rect 22277 9618 22343 9621
rect 27705 9618 27771 9621
rect 22277 9616 27771 9618
rect 22277 9560 22282 9616
rect 22338 9560 27710 9616
rect 27766 9560 27771 9616
rect 22277 9558 27771 9560
rect 22277 9555 22343 9558
rect 27705 9555 27771 9558
rect 17125 9482 17191 9485
rect 21173 9482 21239 9485
rect 24761 9482 24827 9485
rect 17125 9480 21239 9482
rect 17125 9424 17130 9480
rect 17186 9424 21178 9480
rect 21234 9424 21239 9480
rect 17125 9422 21239 9424
rect 17125 9419 17191 9422
rect 21173 9419 21239 9422
rect 21636 9480 24827 9482
rect 21636 9424 24766 9480
rect 24822 9424 24827 9480
rect 21636 9422 24827 9424
rect 19793 9346 19859 9349
rect 21636 9346 21696 9422
rect 24761 9419 24827 9422
rect 19793 9344 21696 9346
rect 19793 9288 19798 9344
rect 19854 9288 21696 9344
rect 19793 9286 21696 9288
rect 21817 9346 21883 9349
rect 24025 9346 24091 9349
rect 21817 9344 24091 9346
rect 21817 9288 21822 9344
rect 21878 9288 24030 9344
rect 24086 9288 24091 9344
rect 21817 9286 24091 9288
rect 19793 9283 19859 9286
rect 21817 9283 21883 9286
rect 24025 9283 24091 9286
rect 14641 9210 14707 9213
rect 17861 9210 17927 9213
rect 14641 9208 17927 9210
rect 14641 9152 14646 9208
rect 14702 9152 17866 9208
rect 17922 9152 17927 9208
rect 14641 9150 17927 9152
rect 14641 9147 14707 9150
rect 17861 9147 17927 9150
rect 20069 9210 20135 9213
rect 24669 9210 24735 9213
rect 20069 9208 24735 9210
rect 20069 9152 20074 9208
rect 20130 9152 24674 9208
rect 24730 9152 24735 9208
rect 20069 9150 24735 9152
rect 20069 9147 20135 9150
rect 24669 9147 24735 9150
rect 12985 9074 13051 9077
rect 17769 9074 17835 9077
rect 12985 9072 17835 9074
rect 12985 9016 12990 9072
rect 13046 9016 17774 9072
rect 17830 9016 17835 9072
rect 12985 9014 17835 9016
rect 12985 9011 13051 9014
rect 17769 9011 17835 9014
rect 21633 9074 21699 9077
rect 22461 9074 22527 9077
rect 21633 9072 22527 9074
rect 21633 9016 21638 9072
rect 21694 9016 22466 9072
rect 22522 9016 22527 9072
rect 21633 9014 22527 9016
rect 21633 9011 21699 9014
rect 22461 9011 22527 9014
rect 13721 8938 13787 8941
rect 28073 8938 28139 8941
rect 13721 8936 28139 8938
rect 13721 8880 13726 8936
rect 13782 8880 28078 8936
rect 28134 8880 28139 8936
rect 13721 8878 28139 8880
rect 13721 8875 13787 8878
rect 28073 8875 28139 8878
rect 21357 8802 21423 8805
rect 22737 8802 22803 8805
rect 21357 8800 22803 8802
rect 21357 8744 21362 8800
rect 21418 8744 22742 8800
rect 22798 8744 22803 8800
rect 21357 8742 22803 8744
rect 21357 8739 21423 8742
rect 22737 8739 22803 8742
rect 12376 8736 12692 8737
rect 12376 8672 12382 8736
rect 12446 8672 12462 8736
rect 12526 8672 12542 8736
rect 12606 8672 12622 8736
rect 12686 8672 12692 8736
rect 12376 8671 12692 8672
rect 23806 8736 24122 8737
rect 23806 8672 23812 8736
rect 23876 8672 23892 8736
rect 23956 8672 23972 8736
rect 24036 8672 24052 8736
rect 24116 8672 24122 8736
rect 23806 8671 24122 8672
rect 35236 8736 35552 8737
rect 35236 8672 35242 8736
rect 35306 8672 35322 8736
rect 35386 8672 35402 8736
rect 35466 8672 35482 8736
rect 35546 8672 35552 8736
rect 35236 8671 35552 8672
rect 46666 8736 46982 8737
rect 46666 8672 46672 8736
rect 46736 8672 46752 8736
rect 46816 8672 46832 8736
rect 46896 8672 46912 8736
rect 46976 8672 46982 8736
rect 46666 8671 46982 8672
rect 19701 8666 19767 8669
rect 22645 8666 22711 8669
rect 19701 8664 22711 8666
rect 19701 8608 19706 8664
rect 19762 8608 22650 8664
rect 22706 8608 22711 8664
rect 19701 8606 22711 8608
rect 19701 8603 19767 8606
rect 22645 8603 22711 8606
rect 14825 8530 14891 8533
rect 25405 8530 25471 8533
rect 14825 8528 25471 8530
rect 14825 8472 14830 8528
rect 14886 8472 25410 8528
rect 25466 8472 25471 8528
rect 14825 8470 25471 8472
rect 14825 8467 14891 8470
rect 25405 8467 25471 8470
rect 14457 8394 14523 8397
rect 20897 8394 20963 8397
rect 14457 8392 20963 8394
rect 14457 8336 14462 8392
rect 14518 8336 20902 8392
rect 20958 8336 20963 8392
rect 14457 8334 20963 8336
rect 14457 8331 14523 8334
rect 20897 8331 20963 8334
rect 21541 8394 21607 8397
rect 23749 8394 23815 8397
rect 21541 8392 23815 8394
rect 21541 8336 21546 8392
rect 21602 8336 23754 8392
rect 23810 8336 23815 8392
rect 21541 8334 23815 8336
rect 21541 8331 21607 8334
rect 23749 8331 23815 8334
rect 24393 8394 24459 8397
rect 28165 8394 28231 8397
rect 24393 8392 28231 8394
rect 24393 8336 24398 8392
rect 24454 8336 28170 8392
rect 28226 8336 28231 8392
rect 24393 8334 28231 8336
rect 24393 8331 24459 8334
rect 28165 8331 28231 8334
rect 11973 8258 12039 8261
rect 16205 8258 16271 8261
rect 11973 8256 16271 8258
rect 11973 8200 11978 8256
rect 12034 8200 16210 8256
rect 16266 8200 16271 8256
rect 11973 8198 16271 8200
rect 11973 8195 12039 8198
rect 16205 8195 16271 8198
rect 19333 8258 19399 8261
rect 21357 8258 21423 8261
rect 19333 8256 21423 8258
rect 19333 8200 19338 8256
rect 19394 8200 21362 8256
rect 21418 8200 21423 8256
rect 19333 8198 21423 8200
rect 19333 8195 19399 8198
rect 21357 8195 21423 8198
rect 23841 8258 23907 8261
rect 28257 8258 28323 8261
rect 23841 8256 28323 8258
rect 23841 8200 23846 8256
rect 23902 8200 28262 8256
rect 28318 8200 28323 8256
rect 23841 8198 28323 8200
rect 23841 8195 23907 8198
rect 28257 8195 28323 8198
rect 6661 8192 6977 8193
rect 6661 8128 6667 8192
rect 6731 8128 6747 8192
rect 6811 8128 6827 8192
rect 6891 8128 6907 8192
rect 6971 8128 6977 8192
rect 6661 8127 6977 8128
rect 18091 8192 18407 8193
rect 18091 8128 18097 8192
rect 18161 8128 18177 8192
rect 18241 8128 18257 8192
rect 18321 8128 18337 8192
rect 18401 8128 18407 8192
rect 18091 8127 18407 8128
rect 29521 8192 29837 8193
rect 29521 8128 29527 8192
rect 29591 8128 29607 8192
rect 29671 8128 29687 8192
rect 29751 8128 29767 8192
rect 29831 8128 29837 8192
rect 29521 8127 29837 8128
rect 40951 8192 41267 8193
rect 40951 8128 40957 8192
rect 41021 8128 41037 8192
rect 41101 8128 41117 8192
rect 41181 8128 41197 8192
rect 41261 8128 41267 8192
rect 40951 8127 41267 8128
rect 18505 8122 18571 8125
rect 35065 8122 35131 8125
rect 18505 8120 26986 8122
rect 18505 8064 18510 8120
rect 18566 8064 26986 8120
rect 18505 8062 26986 8064
rect 18505 8059 18571 8062
rect 17953 7986 18019 7989
rect 26926 7986 26986 8062
rect 30054 8120 35131 8122
rect 30054 8064 35070 8120
rect 35126 8064 35131 8120
rect 30054 8062 35131 8064
rect 30054 7986 30114 8062
rect 35065 8059 35131 8062
rect 35801 7986 35867 7989
rect 17953 7984 26802 7986
rect 17953 7928 17958 7984
rect 18014 7928 26802 7984
rect 17953 7926 26802 7928
rect 26926 7926 30114 7986
rect 31710 7984 35867 7986
rect 31710 7928 35806 7984
rect 35862 7928 35867 7984
rect 31710 7926 35867 7928
rect 17953 7923 18019 7926
rect 2313 7850 2379 7853
rect 26742 7850 26802 7926
rect 31710 7850 31770 7926
rect 35801 7923 35867 7926
rect 2313 7848 24410 7850
rect 2313 7792 2318 7848
rect 2374 7792 24410 7848
rect 2313 7790 24410 7792
rect 26742 7790 31770 7850
rect 2313 7787 2379 7790
rect 15101 7714 15167 7717
rect 19333 7714 19399 7717
rect 15101 7712 19399 7714
rect 15101 7656 15106 7712
rect 15162 7656 19338 7712
rect 19394 7656 19399 7712
rect 15101 7654 19399 7656
rect 15101 7651 15167 7654
rect 19333 7651 19399 7654
rect 22829 7714 22895 7717
rect 24350 7714 24410 7790
rect 26785 7714 26851 7717
rect 22829 7712 23674 7714
rect 22829 7656 22834 7712
rect 22890 7656 23674 7712
rect 22829 7654 23674 7656
rect 24350 7712 26851 7714
rect 24350 7656 26790 7712
rect 26846 7656 26851 7712
rect 24350 7654 26851 7656
rect 22829 7651 22895 7654
rect 12376 7648 12692 7649
rect 12376 7584 12382 7648
rect 12446 7584 12462 7648
rect 12526 7584 12542 7648
rect 12606 7584 12622 7648
rect 12686 7584 12692 7648
rect 12376 7583 12692 7584
rect 14641 7578 14707 7581
rect 16941 7578 17007 7581
rect 14641 7576 17007 7578
rect 14641 7520 14646 7576
rect 14702 7520 16946 7576
rect 17002 7520 17007 7576
rect 14641 7518 17007 7520
rect 14641 7515 14707 7518
rect 16941 7515 17007 7518
rect 18137 7578 18203 7581
rect 21541 7578 21607 7581
rect 18137 7576 21607 7578
rect 18137 7520 18142 7576
rect 18198 7520 21546 7576
rect 21602 7520 21607 7576
rect 18137 7518 21607 7520
rect 18137 7515 18203 7518
rect 21541 7515 21607 7518
rect 16665 7442 16731 7445
rect 23381 7442 23447 7445
rect 16665 7440 23447 7442
rect 16665 7384 16670 7440
rect 16726 7384 23386 7440
rect 23442 7384 23447 7440
rect 16665 7382 23447 7384
rect 23614 7442 23674 7654
rect 26785 7651 26851 7654
rect 23806 7648 24122 7649
rect 23806 7584 23812 7648
rect 23876 7584 23892 7648
rect 23956 7584 23972 7648
rect 24036 7584 24052 7648
rect 24116 7584 24122 7648
rect 23806 7583 24122 7584
rect 35236 7648 35552 7649
rect 35236 7584 35242 7648
rect 35306 7584 35322 7648
rect 35386 7584 35402 7648
rect 35466 7584 35482 7648
rect 35546 7584 35552 7648
rect 35236 7583 35552 7584
rect 46666 7648 46982 7649
rect 46666 7584 46672 7648
rect 46736 7584 46752 7648
rect 46816 7584 46832 7648
rect 46896 7584 46912 7648
rect 46976 7584 46982 7648
rect 46666 7583 46982 7584
rect 38745 7442 38811 7445
rect 23614 7440 38811 7442
rect 23614 7384 38750 7440
rect 38806 7384 38811 7440
rect 23614 7382 38811 7384
rect 16665 7379 16731 7382
rect 23381 7379 23447 7382
rect 38745 7379 38811 7382
rect 14825 7306 14891 7309
rect 29177 7306 29243 7309
rect 14825 7304 29243 7306
rect 14825 7248 14830 7304
rect 14886 7248 29182 7304
rect 29238 7248 29243 7304
rect 14825 7246 29243 7248
rect 14825 7243 14891 7246
rect 29177 7243 29243 7246
rect 19977 7170 20043 7173
rect 27981 7170 28047 7173
rect 19977 7168 28047 7170
rect 19977 7112 19982 7168
rect 20038 7112 27986 7168
rect 28042 7112 28047 7168
rect 19977 7110 28047 7112
rect 19977 7107 20043 7110
rect 27981 7107 28047 7110
rect 6661 7104 6977 7105
rect 6661 7040 6667 7104
rect 6731 7040 6747 7104
rect 6811 7040 6827 7104
rect 6891 7040 6907 7104
rect 6971 7040 6977 7104
rect 6661 7039 6977 7040
rect 18091 7104 18407 7105
rect 18091 7040 18097 7104
rect 18161 7040 18177 7104
rect 18241 7040 18257 7104
rect 18321 7040 18337 7104
rect 18401 7040 18407 7104
rect 18091 7039 18407 7040
rect 29521 7104 29837 7105
rect 29521 7040 29527 7104
rect 29591 7040 29607 7104
rect 29671 7040 29687 7104
rect 29751 7040 29767 7104
rect 29831 7040 29837 7104
rect 29521 7039 29837 7040
rect 40951 7104 41267 7105
rect 40951 7040 40957 7104
rect 41021 7040 41037 7104
rect 41101 7040 41117 7104
rect 41181 7040 41197 7104
rect 41261 7040 41267 7104
rect 40951 7039 41267 7040
rect 3233 6898 3299 6901
rect 26233 6898 26299 6901
rect 3233 6896 26299 6898
rect 3233 6840 3238 6896
rect 3294 6840 26238 6896
rect 26294 6840 26299 6896
rect 3233 6838 26299 6840
rect 3233 6835 3299 6838
rect 26233 6835 26299 6838
rect 12376 6560 12692 6561
rect 12376 6496 12382 6560
rect 12446 6496 12462 6560
rect 12526 6496 12542 6560
rect 12606 6496 12622 6560
rect 12686 6496 12692 6560
rect 12376 6495 12692 6496
rect 23806 6560 24122 6561
rect 23806 6496 23812 6560
rect 23876 6496 23892 6560
rect 23956 6496 23972 6560
rect 24036 6496 24052 6560
rect 24116 6496 24122 6560
rect 23806 6495 24122 6496
rect 35236 6560 35552 6561
rect 35236 6496 35242 6560
rect 35306 6496 35322 6560
rect 35386 6496 35402 6560
rect 35466 6496 35482 6560
rect 35546 6496 35552 6560
rect 35236 6495 35552 6496
rect 46666 6560 46982 6561
rect 46666 6496 46672 6560
rect 46736 6496 46752 6560
rect 46816 6496 46832 6560
rect 46896 6496 46912 6560
rect 46976 6496 46982 6560
rect 46666 6495 46982 6496
rect 6661 6016 6977 6017
rect 6661 5952 6667 6016
rect 6731 5952 6747 6016
rect 6811 5952 6827 6016
rect 6891 5952 6907 6016
rect 6971 5952 6977 6016
rect 6661 5951 6977 5952
rect 18091 6016 18407 6017
rect 18091 5952 18097 6016
rect 18161 5952 18177 6016
rect 18241 5952 18257 6016
rect 18321 5952 18337 6016
rect 18401 5952 18407 6016
rect 18091 5951 18407 5952
rect 29521 6016 29837 6017
rect 29521 5952 29527 6016
rect 29591 5952 29607 6016
rect 29671 5952 29687 6016
rect 29751 5952 29767 6016
rect 29831 5952 29837 6016
rect 29521 5951 29837 5952
rect 40951 6016 41267 6017
rect 40951 5952 40957 6016
rect 41021 5952 41037 6016
rect 41101 5952 41117 6016
rect 41181 5952 41197 6016
rect 41261 5952 41267 6016
rect 40951 5951 41267 5952
rect 12376 5472 12692 5473
rect 12376 5408 12382 5472
rect 12446 5408 12462 5472
rect 12526 5408 12542 5472
rect 12606 5408 12622 5472
rect 12686 5408 12692 5472
rect 12376 5407 12692 5408
rect 23806 5472 24122 5473
rect 23806 5408 23812 5472
rect 23876 5408 23892 5472
rect 23956 5408 23972 5472
rect 24036 5408 24052 5472
rect 24116 5408 24122 5472
rect 23806 5407 24122 5408
rect 35236 5472 35552 5473
rect 35236 5408 35242 5472
rect 35306 5408 35322 5472
rect 35386 5408 35402 5472
rect 35466 5408 35482 5472
rect 35546 5408 35552 5472
rect 35236 5407 35552 5408
rect 46666 5472 46982 5473
rect 46666 5408 46672 5472
rect 46736 5408 46752 5472
rect 46816 5408 46832 5472
rect 46896 5408 46912 5472
rect 46976 5408 46982 5472
rect 46666 5407 46982 5408
rect 6661 4928 6977 4929
rect 6661 4864 6667 4928
rect 6731 4864 6747 4928
rect 6811 4864 6827 4928
rect 6891 4864 6907 4928
rect 6971 4864 6977 4928
rect 6661 4863 6977 4864
rect 18091 4928 18407 4929
rect 18091 4864 18097 4928
rect 18161 4864 18177 4928
rect 18241 4864 18257 4928
rect 18321 4864 18337 4928
rect 18401 4864 18407 4928
rect 18091 4863 18407 4864
rect 29521 4928 29837 4929
rect 29521 4864 29527 4928
rect 29591 4864 29607 4928
rect 29671 4864 29687 4928
rect 29751 4864 29767 4928
rect 29831 4864 29837 4928
rect 29521 4863 29837 4864
rect 40951 4928 41267 4929
rect 40951 4864 40957 4928
rect 41021 4864 41037 4928
rect 41101 4864 41117 4928
rect 41181 4864 41197 4928
rect 41261 4864 41267 4928
rect 40951 4863 41267 4864
rect 12376 4384 12692 4385
rect 12376 4320 12382 4384
rect 12446 4320 12462 4384
rect 12526 4320 12542 4384
rect 12606 4320 12622 4384
rect 12686 4320 12692 4384
rect 12376 4319 12692 4320
rect 23806 4384 24122 4385
rect 23806 4320 23812 4384
rect 23876 4320 23892 4384
rect 23956 4320 23972 4384
rect 24036 4320 24052 4384
rect 24116 4320 24122 4384
rect 23806 4319 24122 4320
rect 35236 4384 35552 4385
rect 35236 4320 35242 4384
rect 35306 4320 35322 4384
rect 35386 4320 35402 4384
rect 35466 4320 35482 4384
rect 35546 4320 35552 4384
rect 35236 4319 35552 4320
rect 46666 4384 46982 4385
rect 46666 4320 46672 4384
rect 46736 4320 46752 4384
rect 46816 4320 46832 4384
rect 46896 4320 46912 4384
rect 46976 4320 46982 4384
rect 46666 4319 46982 4320
rect 6661 3840 6977 3841
rect 6661 3776 6667 3840
rect 6731 3776 6747 3840
rect 6811 3776 6827 3840
rect 6891 3776 6907 3840
rect 6971 3776 6977 3840
rect 6661 3775 6977 3776
rect 18091 3840 18407 3841
rect 18091 3776 18097 3840
rect 18161 3776 18177 3840
rect 18241 3776 18257 3840
rect 18321 3776 18337 3840
rect 18401 3776 18407 3840
rect 18091 3775 18407 3776
rect 29521 3840 29837 3841
rect 29521 3776 29527 3840
rect 29591 3776 29607 3840
rect 29671 3776 29687 3840
rect 29751 3776 29767 3840
rect 29831 3776 29837 3840
rect 29521 3775 29837 3776
rect 40951 3840 41267 3841
rect 40951 3776 40957 3840
rect 41021 3776 41037 3840
rect 41101 3776 41117 3840
rect 41181 3776 41197 3840
rect 41261 3776 41267 3840
rect 40951 3775 41267 3776
rect 12376 3296 12692 3297
rect 12376 3232 12382 3296
rect 12446 3232 12462 3296
rect 12526 3232 12542 3296
rect 12606 3232 12622 3296
rect 12686 3232 12692 3296
rect 12376 3231 12692 3232
rect 23806 3296 24122 3297
rect 23806 3232 23812 3296
rect 23876 3232 23892 3296
rect 23956 3232 23972 3296
rect 24036 3232 24052 3296
rect 24116 3232 24122 3296
rect 23806 3231 24122 3232
rect 35236 3296 35552 3297
rect 35236 3232 35242 3296
rect 35306 3232 35322 3296
rect 35386 3232 35402 3296
rect 35466 3232 35482 3296
rect 35546 3232 35552 3296
rect 35236 3231 35552 3232
rect 46666 3296 46982 3297
rect 46666 3232 46672 3296
rect 46736 3232 46752 3296
rect 46816 3232 46832 3296
rect 46896 3232 46912 3296
rect 46976 3232 46982 3296
rect 46666 3231 46982 3232
rect 6661 2752 6977 2753
rect 6661 2688 6667 2752
rect 6731 2688 6747 2752
rect 6811 2688 6827 2752
rect 6891 2688 6907 2752
rect 6971 2688 6977 2752
rect 6661 2687 6977 2688
rect 18091 2752 18407 2753
rect 18091 2688 18097 2752
rect 18161 2688 18177 2752
rect 18241 2688 18257 2752
rect 18321 2688 18337 2752
rect 18401 2688 18407 2752
rect 18091 2687 18407 2688
rect 29521 2752 29837 2753
rect 29521 2688 29527 2752
rect 29591 2688 29607 2752
rect 29671 2688 29687 2752
rect 29751 2688 29767 2752
rect 29831 2688 29837 2752
rect 29521 2687 29837 2688
rect 40951 2752 41267 2753
rect 40951 2688 40957 2752
rect 41021 2688 41037 2752
rect 41101 2688 41117 2752
rect 41181 2688 41197 2752
rect 41261 2688 41267 2752
rect 40951 2687 41267 2688
rect 12376 2208 12692 2209
rect 12376 2144 12382 2208
rect 12446 2144 12462 2208
rect 12526 2144 12542 2208
rect 12606 2144 12622 2208
rect 12686 2144 12692 2208
rect 12376 2143 12692 2144
rect 23806 2208 24122 2209
rect 23806 2144 23812 2208
rect 23876 2144 23892 2208
rect 23956 2144 23972 2208
rect 24036 2144 24052 2208
rect 24116 2144 24122 2208
rect 23806 2143 24122 2144
rect 35236 2208 35552 2209
rect 35236 2144 35242 2208
rect 35306 2144 35322 2208
rect 35386 2144 35402 2208
rect 35466 2144 35482 2208
rect 35546 2144 35552 2208
rect 35236 2143 35552 2144
rect 46666 2208 46982 2209
rect 46666 2144 46672 2208
rect 46736 2144 46752 2208
rect 46816 2144 46832 2208
rect 46896 2144 46912 2208
rect 46976 2144 46982 2208
rect 46666 2143 46982 2144
rect 6661 1664 6977 1665
rect 6661 1600 6667 1664
rect 6731 1600 6747 1664
rect 6811 1600 6827 1664
rect 6891 1600 6907 1664
rect 6971 1600 6977 1664
rect 6661 1599 6977 1600
rect 18091 1664 18407 1665
rect 18091 1600 18097 1664
rect 18161 1600 18177 1664
rect 18241 1600 18257 1664
rect 18321 1600 18337 1664
rect 18401 1600 18407 1664
rect 18091 1599 18407 1600
rect 29521 1664 29837 1665
rect 29521 1600 29527 1664
rect 29591 1600 29607 1664
rect 29671 1600 29687 1664
rect 29751 1600 29767 1664
rect 29831 1600 29837 1664
rect 29521 1599 29837 1600
rect 40951 1664 41267 1665
rect 40951 1600 40957 1664
rect 41021 1600 41037 1664
rect 41101 1600 41117 1664
rect 41181 1600 41197 1664
rect 41261 1600 41267 1664
rect 40951 1599 41267 1600
rect 12376 1120 12692 1121
rect 12376 1056 12382 1120
rect 12446 1056 12462 1120
rect 12526 1056 12542 1120
rect 12606 1056 12622 1120
rect 12686 1056 12692 1120
rect 12376 1055 12692 1056
rect 23806 1120 24122 1121
rect 23806 1056 23812 1120
rect 23876 1056 23892 1120
rect 23956 1056 23972 1120
rect 24036 1056 24052 1120
rect 24116 1056 24122 1120
rect 23806 1055 24122 1056
rect 35236 1120 35552 1121
rect 35236 1056 35242 1120
rect 35306 1056 35322 1120
rect 35386 1056 35402 1120
rect 35466 1056 35482 1120
rect 35546 1056 35552 1120
rect 35236 1055 35552 1056
rect 46666 1120 46982 1121
rect 46666 1056 46672 1120
rect 46736 1056 46752 1120
rect 46816 1056 46832 1120
rect 46896 1056 46912 1120
rect 46976 1056 46982 1120
rect 46666 1055 46982 1056
<< via3 >>
rect 12382 8732 12446 8736
rect 12382 8676 12386 8732
rect 12386 8676 12442 8732
rect 12442 8676 12446 8732
rect 12382 8672 12446 8676
rect 12462 8732 12526 8736
rect 12462 8676 12466 8732
rect 12466 8676 12522 8732
rect 12522 8676 12526 8732
rect 12462 8672 12526 8676
rect 12542 8732 12606 8736
rect 12542 8676 12546 8732
rect 12546 8676 12602 8732
rect 12602 8676 12606 8732
rect 12542 8672 12606 8676
rect 12622 8732 12686 8736
rect 12622 8676 12626 8732
rect 12626 8676 12682 8732
rect 12682 8676 12686 8732
rect 12622 8672 12686 8676
rect 23812 8732 23876 8736
rect 23812 8676 23816 8732
rect 23816 8676 23872 8732
rect 23872 8676 23876 8732
rect 23812 8672 23876 8676
rect 23892 8732 23956 8736
rect 23892 8676 23896 8732
rect 23896 8676 23952 8732
rect 23952 8676 23956 8732
rect 23892 8672 23956 8676
rect 23972 8732 24036 8736
rect 23972 8676 23976 8732
rect 23976 8676 24032 8732
rect 24032 8676 24036 8732
rect 23972 8672 24036 8676
rect 24052 8732 24116 8736
rect 24052 8676 24056 8732
rect 24056 8676 24112 8732
rect 24112 8676 24116 8732
rect 24052 8672 24116 8676
rect 35242 8732 35306 8736
rect 35242 8676 35246 8732
rect 35246 8676 35302 8732
rect 35302 8676 35306 8732
rect 35242 8672 35306 8676
rect 35322 8732 35386 8736
rect 35322 8676 35326 8732
rect 35326 8676 35382 8732
rect 35382 8676 35386 8732
rect 35322 8672 35386 8676
rect 35402 8732 35466 8736
rect 35402 8676 35406 8732
rect 35406 8676 35462 8732
rect 35462 8676 35466 8732
rect 35402 8672 35466 8676
rect 35482 8732 35546 8736
rect 35482 8676 35486 8732
rect 35486 8676 35542 8732
rect 35542 8676 35546 8732
rect 35482 8672 35546 8676
rect 46672 8732 46736 8736
rect 46672 8676 46676 8732
rect 46676 8676 46732 8732
rect 46732 8676 46736 8732
rect 46672 8672 46736 8676
rect 46752 8732 46816 8736
rect 46752 8676 46756 8732
rect 46756 8676 46812 8732
rect 46812 8676 46816 8732
rect 46752 8672 46816 8676
rect 46832 8732 46896 8736
rect 46832 8676 46836 8732
rect 46836 8676 46892 8732
rect 46892 8676 46896 8732
rect 46832 8672 46896 8676
rect 46912 8732 46976 8736
rect 46912 8676 46916 8732
rect 46916 8676 46972 8732
rect 46972 8676 46976 8732
rect 46912 8672 46976 8676
rect 6667 8188 6731 8192
rect 6667 8132 6671 8188
rect 6671 8132 6727 8188
rect 6727 8132 6731 8188
rect 6667 8128 6731 8132
rect 6747 8188 6811 8192
rect 6747 8132 6751 8188
rect 6751 8132 6807 8188
rect 6807 8132 6811 8188
rect 6747 8128 6811 8132
rect 6827 8188 6891 8192
rect 6827 8132 6831 8188
rect 6831 8132 6887 8188
rect 6887 8132 6891 8188
rect 6827 8128 6891 8132
rect 6907 8188 6971 8192
rect 6907 8132 6911 8188
rect 6911 8132 6967 8188
rect 6967 8132 6971 8188
rect 6907 8128 6971 8132
rect 18097 8188 18161 8192
rect 18097 8132 18101 8188
rect 18101 8132 18157 8188
rect 18157 8132 18161 8188
rect 18097 8128 18161 8132
rect 18177 8188 18241 8192
rect 18177 8132 18181 8188
rect 18181 8132 18237 8188
rect 18237 8132 18241 8188
rect 18177 8128 18241 8132
rect 18257 8188 18321 8192
rect 18257 8132 18261 8188
rect 18261 8132 18317 8188
rect 18317 8132 18321 8188
rect 18257 8128 18321 8132
rect 18337 8188 18401 8192
rect 18337 8132 18341 8188
rect 18341 8132 18397 8188
rect 18397 8132 18401 8188
rect 18337 8128 18401 8132
rect 29527 8188 29591 8192
rect 29527 8132 29531 8188
rect 29531 8132 29587 8188
rect 29587 8132 29591 8188
rect 29527 8128 29591 8132
rect 29607 8188 29671 8192
rect 29607 8132 29611 8188
rect 29611 8132 29667 8188
rect 29667 8132 29671 8188
rect 29607 8128 29671 8132
rect 29687 8188 29751 8192
rect 29687 8132 29691 8188
rect 29691 8132 29747 8188
rect 29747 8132 29751 8188
rect 29687 8128 29751 8132
rect 29767 8188 29831 8192
rect 29767 8132 29771 8188
rect 29771 8132 29827 8188
rect 29827 8132 29831 8188
rect 29767 8128 29831 8132
rect 40957 8188 41021 8192
rect 40957 8132 40961 8188
rect 40961 8132 41017 8188
rect 41017 8132 41021 8188
rect 40957 8128 41021 8132
rect 41037 8188 41101 8192
rect 41037 8132 41041 8188
rect 41041 8132 41097 8188
rect 41097 8132 41101 8188
rect 41037 8128 41101 8132
rect 41117 8188 41181 8192
rect 41117 8132 41121 8188
rect 41121 8132 41177 8188
rect 41177 8132 41181 8188
rect 41117 8128 41181 8132
rect 41197 8188 41261 8192
rect 41197 8132 41201 8188
rect 41201 8132 41257 8188
rect 41257 8132 41261 8188
rect 41197 8128 41261 8132
rect 12382 7644 12446 7648
rect 12382 7588 12386 7644
rect 12386 7588 12442 7644
rect 12442 7588 12446 7644
rect 12382 7584 12446 7588
rect 12462 7644 12526 7648
rect 12462 7588 12466 7644
rect 12466 7588 12522 7644
rect 12522 7588 12526 7644
rect 12462 7584 12526 7588
rect 12542 7644 12606 7648
rect 12542 7588 12546 7644
rect 12546 7588 12602 7644
rect 12602 7588 12606 7644
rect 12542 7584 12606 7588
rect 12622 7644 12686 7648
rect 12622 7588 12626 7644
rect 12626 7588 12682 7644
rect 12682 7588 12686 7644
rect 12622 7584 12686 7588
rect 23812 7644 23876 7648
rect 23812 7588 23816 7644
rect 23816 7588 23872 7644
rect 23872 7588 23876 7644
rect 23812 7584 23876 7588
rect 23892 7644 23956 7648
rect 23892 7588 23896 7644
rect 23896 7588 23952 7644
rect 23952 7588 23956 7644
rect 23892 7584 23956 7588
rect 23972 7644 24036 7648
rect 23972 7588 23976 7644
rect 23976 7588 24032 7644
rect 24032 7588 24036 7644
rect 23972 7584 24036 7588
rect 24052 7644 24116 7648
rect 24052 7588 24056 7644
rect 24056 7588 24112 7644
rect 24112 7588 24116 7644
rect 24052 7584 24116 7588
rect 35242 7644 35306 7648
rect 35242 7588 35246 7644
rect 35246 7588 35302 7644
rect 35302 7588 35306 7644
rect 35242 7584 35306 7588
rect 35322 7644 35386 7648
rect 35322 7588 35326 7644
rect 35326 7588 35382 7644
rect 35382 7588 35386 7644
rect 35322 7584 35386 7588
rect 35402 7644 35466 7648
rect 35402 7588 35406 7644
rect 35406 7588 35462 7644
rect 35462 7588 35466 7644
rect 35402 7584 35466 7588
rect 35482 7644 35546 7648
rect 35482 7588 35486 7644
rect 35486 7588 35542 7644
rect 35542 7588 35546 7644
rect 35482 7584 35546 7588
rect 46672 7644 46736 7648
rect 46672 7588 46676 7644
rect 46676 7588 46732 7644
rect 46732 7588 46736 7644
rect 46672 7584 46736 7588
rect 46752 7644 46816 7648
rect 46752 7588 46756 7644
rect 46756 7588 46812 7644
rect 46812 7588 46816 7644
rect 46752 7584 46816 7588
rect 46832 7644 46896 7648
rect 46832 7588 46836 7644
rect 46836 7588 46892 7644
rect 46892 7588 46896 7644
rect 46832 7584 46896 7588
rect 46912 7644 46976 7648
rect 46912 7588 46916 7644
rect 46916 7588 46972 7644
rect 46972 7588 46976 7644
rect 46912 7584 46976 7588
rect 6667 7100 6731 7104
rect 6667 7044 6671 7100
rect 6671 7044 6727 7100
rect 6727 7044 6731 7100
rect 6667 7040 6731 7044
rect 6747 7100 6811 7104
rect 6747 7044 6751 7100
rect 6751 7044 6807 7100
rect 6807 7044 6811 7100
rect 6747 7040 6811 7044
rect 6827 7100 6891 7104
rect 6827 7044 6831 7100
rect 6831 7044 6887 7100
rect 6887 7044 6891 7100
rect 6827 7040 6891 7044
rect 6907 7100 6971 7104
rect 6907 7044 6911 7100
rect 6911 7044 6967 7100
rect 6967 7044 6971 7100
rect 6907 7040 6971 7044
rect 18097 7100 18161 7104
rect 18097 7044 18101 7100
rect 18101 7044 18157 7100
rect 18157 7044 18161 7100
rect 18097 7040 18161 7044
rect 18177 7100 18241 7104
rect 18177 7044 18181 7100
rect 18181 7044 18237 7100
rect 18237 7044 18241 7100
rect 18177 7040 18241 7044
rect 18257 7100 18321 7104
rect 18257 7044 18261 7100
rect 18261 7044 18317 7100
rect 18317 7044 18321 7100
rect 18257 7040 18321 7044
rect 18337 7100 18401 7104
rect 18337 7044 18341 7100
rect 18341 7044 18397 7100
rect 18397 7044 18401 7100
rect 18337 7040 18401 7044
rect 29527 7100 29591 7104
rect 29527 7044 29531 7100
rect 29531 7044 29587 7100
rect 29587 7044 29591 7100
rect 29527 7040 29591 7044
rect 29607 7100 29671 7104
rect 29607 7044 29611 7100
rect 29611 7044 29667 7100
rect 29667 7044 29671 7100
rect 29607 7040 29671 7044
rect 29687 7100 29751 7104
rect 29687 7044 29691 7100
rect 29691 7044 29747 7100
rect 29747 7044 29751 7100
rect 29687 7040 29751 7044
rect 29767 7100 29831 7104
rect 29767 7044 29771 7100
rect 29771 7044 29827 7100
rect 29827 7044 29831 7100
rect 29767 7040 29831 7044
rect 40957 7100 41021 7104
rect 40957 7044 40961 7100
rect 40961 7044 41017 7100
rect 41017 7044 41021 7100
rect 40957 7040 41021 7044
rect 41037 7100 41101 7104
rect 41037 7044 41041 7100
rect 41041 7044 41097 7100
rect 41097 7044 41101 7100
rect 41037 7040 41101 7044
rect 41117 7100 41181 7104
rect 41117 7044 41121 7100
rect 41121 7044 41177 7100
rect 41177 7044 41181 7100
rect 41117 7040 41181 7044
rect 41197 7100 41261 7104
rect 41197 7044 41201 7100
rect 41201 7044 41257 7100
rect 41257 7044 41261 7100
rect 41197 7040 41261 7044
rect 12382 6556 12446 6560
rect 12382 6500 12386 6556
rect 12386 6500 12442 6556
rect 12442 6500 12446 6556
rect 12382 6496 12446 6500
rect 12462 6556 12526 6560
rect 12462 6500 12466 6556
rect 12466 6500 12522 6556
rect 12522 6500 12526 6556
rect 12462 6496 12526 6500
rect 12542 6556 12606 6560
rect 12542 6500 12546 6556
rect 12546 6500 12602 6556
rect 12602 6500 12606 6556
rect 12542 6496 12606 6500
rect 12622 6556 12686 6560
rect 12622 6500 12626 6556
rect 12626 6500 12682 6556
rect 12682 6500 12686 6556
rect 12622 6496 12686 6500
rect 23812 6556 23876 6560
rect 23812 6500 23816 6556
rect 23816 6500 23872 6556
rect 23872 6500 23876 6556
rect 23812 6496 23876 6500
rect 23892 6556 23956 6560
rect 23892 6500 23896 6556
rect 23896 6500 23952 6556
rect 23952 6500 23956 6556
rect 23892 6496 23956 6500
rect 23972 6556 24036 6560
rect 23972 6500 23976 6556
rect 23976 6500 24032 6556
rect 24032 6500 24036 6556
rect 23972 6496 24036 6500
rect 24052 6556 24116 6560
rect 24052 6500 24056 6556
rect 24056 6500 24112 6556
rect 24112 6500 24116 6556
rect 24052 6496 24116 6500
rect 35242 6556 35306 6560
rect 35242 6500 35246 6556
rect 35246 6500 35302 6556
rect 35302 6500 35306 6556
rect 35242 6496 35306 6500
rect 35322 6556 35386 6560
rect 35322 6500 35326 6556
rect 35326 6500 35382 6556
rect 35382 6500 35386 6556
rect 35322 6496 35386 6500
rect 35402 6556 35466 6560
rect 35402 6500 35406 6556
rect 35406 6500 35462 6556
rect 35462 6500 35466 6556
rect 35402 6496 35466 6500
rect 35482 6556 35546 6560
rect 35482 6500 35486 6556
rect 35486 6500 35542 6556
rect 35542 6500 35546 6556
rect 35482 6496 35546 6500
rect 46672 6556 46736 6560
rect 46672 6500 46676 6556
rect 46676 6500 46732 6556
rect 46732 6500 46736 6556
rect 46672 6496 46736 6500
rect 46752 6556 46816 6560
rect 46752 6500 46756 6556
rect 46756 6500 46812 6556
rect 46812 6500 46816 6556
rect 46752 6496 46816 6500
rect 46832 6556 46896 6560
rect 46832 6500 46836 6556
rect 46836 6500 46892 6556
rect 46892 6500 46896 6556
rect 46832 6496 46896 6500
rect 46912 6556 46976 6560
rect 46912 6500 46916 6556
rect 46916 6500 46972 6556
rect 46972 6500 46976 6556
rect 46912 6496 46976 6500
rect 6667 6012 6731 6016
rect 6667 5956 6671 6012
rect 6671 5956 6727 6012
rect 6727 5956 6731 6012
rect 6667 5952 6731 5956
rect 6747 6012 6811 6016
rect 6747 5956 6751 6012
rect 6751 5956 6807 6012
rect 6807 5956 6811 6012
rect 6747 5952 6811 5956
rect 6827 6012 6891 6016
rect 6827 5956 6831 6012
rect 6831 5956 6887 6012
rect 6887 5956 6891 6012
rect 6827 5952 6891 5956
rect 6907 6012 6971 6016
rect 6907 5956 6911 6012
rect 6911 5956 6967 6012
rect 6967 5956 6971 6012
rect 6907 5952 6971 5956
rect 18097 6012 18161 6016
rect 18097 5956 18101 6012
rect 18101 5956 18157 6012
rect 18157 5956 18161 6012
rect 18097 5952 18161 5956
rect 18177 6012 18241 6016
rect 18177 5956 18181 6012
rect 18181 5956 18237 6012
rect 18237 5956 18241 6012
rect 18177 5952 18241 5956
rect 18257 6012 18321 6016
rect 18257 5956 18261 6012
rect 18261 5956 18317 6012
rect 18317 5956 18321 6012
rect 18257 5952 18321 5956
rect 18337 6012 18401 6016
rect 18337 5956 18341 6012
rect 18341 5956 18397 6012
rect 18397 5956 18401 6012
rect 18337 5952 18401 5956
rect 29527 6012 29591 6016
rect 29527 5956 29531 6012
rect 29531 5956 29587 6012
rect 29587 5956 29591 6012
rect 29527 5952 29591 5956
rect 29607 6012 29671 6016
rect 29607 5956 29611 6012
rect 29611 5956 29667 6012
rect 29667 5956 29671 6012
rect 29607 5952 29671 5956
rect 29687 6012 29751 6016
rect 29687 5956 29691 6012
rect 29691 5956 29747 6012
rect 29747 5956 29751 6012
rect 29687 5952 29751 5956
rect 29767 6012 29831 6016
rect 29767 5956 29771 6012
rect 29771 5956 29827 6012
rect 29827 5956 29831 6012
rect 29767 5952 29831 5956
rect 40957 6012 41021 6016
rect 40957 5956 40961 6012
rect 40961 5956 41017 6012
rect 41017 5956 41021 6012
rect 40957 5952 41021 5956
rect 41037 6012 41101 6016
rect 41037 5956 41041 6012
rect 41041 5956 41097 6012
rect 41097 5956 41101 6012
rect 41037 5952 41101 5956
rect 41117 6012 41181 6016
rect 41117 5956 41121 6012
rect 41121 5956 41177 6012
rect 41177 5956 41181 6012
rect 41117 5952 41181 5956
rect 41197 6012 41261 6016
rect 41197 5956 41201 6012
rect 41201 5956 41257 6012
rect 41257 5956 41261 6012
rect 41197 5952 41261 5956
rect 12382 5468 12446 5472
rect 12382 5412 12386 5468
rect 12386 5412 12442 5468
rect 12442 5412 12446 5468
rect 12382 5408 12446 5412
rect 12462 5468 12526 5472
rect 12462 5412 12466 5468
rect 12466 5412 12522 5468
rect 12522 5412 12526 5468
rect 12462 5408 12526 5412
rect 12542 5468 12606 5472
rect 12542 5412 12546 5468
rect 12546 5412 12602 5468
rect 12602 5412 12606 5468
rect 12542 5408 12606 5412
rect 12622 5468 12686 5472
rect 12622 5412 12626 5468
rect 12626 5412 12682 5468
rect 12682 5412 12686 5468
rect 12622 5408 12686 5412
rect 23812 5468 23876 5472
rect 23812 5412 23816 5468
rect 23816 5412 23872 5468
rect 23872 5412 23876 5468
rect 23812 5408 23876 5412
rect 23892 5468 23956 5472
rect 23892 5412 23896 5468
rect 23896 5412 23952 5468
rect 23952 5412 23956 5468
rect 23892 5408 23956 5412
rect 23972 5468 24036 5472
rect 23972 5412 23976 5468
rect 23976 5412 24032 5468
rect 24032 5412 24036 5468
rect 23972 5408 24036 5412
rect 24052 5468 24116 5472
rect 24052 5412 24056 5468
rect 24056 5412 24112 5468
rect 24112 5412 24116 5468
rect 24052 5408 24116 5412
rect 35242 5468 35306 5472
rect 35242 5412 35246 5468
rect 35246 5412 35302 5468
rect 35302 5412 35306 5468
rect 35242 5408 35306 5412
rect 35322 5468 35386 5472
rect 35322 5412 35326 5468
rect 35326 5412 35382 5468
rect 35382 5412 35386 5468
rect 35322 5408 35386 5412
rect 35402 5468 35466 5472
rect 35402 5412 35406 5468
rect 35406 5412 35462 5468
rect 35462 5412 35466 5468
rect 35402 5408 35466 5412
rect 35482 5468 35546 5472
rect 35482 5412 35486 5468
rect 35486 5412 35542 5468
rect 35542 5412 35546 5468
rect 35482 5408 35546 5412
rect 46672 5468 46736 5472
rect 46672 5412 46676 5468
rect 46676 5412 46732 5468
rect 46732 5412 46736 5468
rect 46672 5408 46736 5412
rect 46752 5468 46816 5472
rect 46752 5412 46756 5468
rect 46756 5412 46812 5468
rect 46812 5412 46816 5468
rect 46752 5408 46816 5412
rect 46832 5468 46896 5472
rect 46832 5412 46836 5468
rect 46836 5412 46892 5468
rect 46892 5412 46896 5468
rect 46832 5408 46896 5412
rect 46912 5468 46976 5472
rect 46912 5412 46916 5468
rect 46916 5412 46972 5468
rect 46972 5412 46976 5468
rect 46912 5408 46976 5412
rect 6667 4924 6731 4928
rect 6667 4868 6671 4924
rect 6671 4868 6727 4924
rect 6727 4868 6731 4924
rect 6667 4864 6731 4868
rect 6747 4924 6811 4928
rect 6747 4868 6751 4924
rect 6751 4868 6807 4924
rect 6807 4868 6811 4924
rect 6747 4864 6811 4868
rect 6827 4924 6891 4928
rect 6827 4868 6831 4924
rect 6831 4868 6887 4924
rect 6887 4868 6891 4924
rect 6827 4864 6891 4868
rect 6907 4924 6971 4928
rect 6907 4868 6911 4924
rect 6911 4868 6967 4924
rect 6967 4868 6971 4924
rect 6907 4864 6971 4868
rect 18097 4924 18161 4928
rect 18097 4868 18101 4924
rect 18101 4868 18157 4924
rect 18157 4868 18161 4924
rect 18097 4864 18161 4868
rect 18177 4924 18241 4928
rect 18177 4868 18181 4924
rect 18181 4868 18237 4924
rect 18237 4868 18241 4924
rect 18177 4864 18241 4868
rect 18257 4924 18321 4928
rect 18257 4868 18261 4924
rect 18261 4868 18317 4924
rect 18317 4868 18321 4924
rect 18257 4864 18321 4868
rect 18337 4924 18401 4928
rect 18337 4868 18341 4924
rect 18341 4868 18397 4924
rect 18397 4868 18401 4924
rect 18337 4864 18401 4868
rect 29527 4924 29591 4928
rect 29527 4868 29531 4924
rect 29531 4868 29587 4924
rect 29587 4868 29591 4924
rect 29527 4864 29591 4868
rect 29607 4924 29671 4928
rect 29607 4868 29611 4924
rect 29611 4868 29667 4924
rect 29667 4868 29671 4924
rect 29607 4864 29671 4868
rect 29687 4924 29751 4928
rect 29687 4868 29691 4924
rect 29691 4868 29747 4924
rect 29747 4868 29751 4924
rect 29687 4864 29751 4868
rect 29767 4924 29831 4928
rect 29767 4868 29771 4924
rect 29771 4868 29827 4924
rect 29827 4868 29831 4924
rect 29767 4864 29831 4868
rect 40957 4924 41021 4928
rect 40957 4868 40961 4924
rect 40961 4868 41017 4924
rect 41017 4868 41021 4924
rect 40957 4864 41021 4868
rect 41037 4924 41101 4928
rect 41037 4868 41041 4924
rect 41041 4868 41097 4924
rect 41097 4868 41101 4924
rect 41037 4864 41101 4868
rect 41117 4924 41181 4928
rect 41117 4868 41121 4924
rect 41121 4868 41177 4924
rect 41177 4868 41181 4924
rect 41117 4864 41181 4868
rect 41197 4924 41261 4928
rect 41197 4868 41201 4924
rect 41201 4868 41257 4924
rect 41257 4868 41261 4924
rect 41197 4864 41261 4868
rect 12382 4380 12446 4384
rect 12382 4324 12386 4380
rect 12386 4324 12442 4380
rect 12442 4324 12446 4380
rect 12382 4320 12446 4324
rect 12462 4380 12526 4384
rect 12462 4324 12466 4380
rect 12466 4324 12522 4380
rect 12522 4324 12526 4380
rect 12462 4320 12526 4324
rect 12542 4380 12606 4384
rect 12542 4324 12546 4380
rect 12546 4324 12602 4380
rect 12602 4324 12606 4380
rect 12542 4320 12606 4324
rect 12622 4380 12686 4384
rect 12622 4324 12626 4380
rect 12626 4324 12682 4380
rect 12682 4324 12686 4380
rect 12622 4320 12686 4324
rect 23812 4380 23876 4384
rect 23812 4324 23816 4380
rect 23816 4324 23872 4380
rect 23872 4324 23876 4380
rect 23812 4320 23876 4324
rect 23892 4380 23956 4384
rect 23892 4324 23896 4380
rect 23896 4324 23952 4380
rect 23952 4324 23956 4380
rect 23892 4320 23956 4324
rect 23972 4380 24036 4384
rect 23972 4324 23976 4380
rect 23976 4324 24032 4380
rect 24032 4324 24036 4380
rect 23972 4320 24036 4324
rect 24052 4380 24116 4384
rect 24052 4324 24056 4380
rect 24056 4324 24112 4380
rect 24112 4324 24116 4380
rect 24052 4320 24116 4324
rect 35242 4380 35306 4384
rect 35242 4324 35246 4380
rect 35246 4324 35302 4380
rect 35302 4324 35306 4380
rect 35242 4320 35306 4324
rect 35322 4380 35386 4384
rect 35322 4324 35326 4380
rect 35326 4324 35382 4380
rect 35382 4324 35386 4380
rect 35322 4320 35386 4324
rect 35402 4380 35466 4384
rect 35402 4324 35406 4380
rect 35406 4324 35462 4380
rect 35462 4324 35466 4380
rect 35402 4320 35466 4324
rect 35482 4380 35546 4384
rect 35482 4324 35486 4380
rect 35486 4324 35542 4380
rect 35542 4324 35546 4380
rect 35482 4320 35546 4324
rect 46672 4380 46736 4384
rect 46672 4324 46676 4380
rect 46676 4324 46732 4380
rect 46732 4324 46736 4380
rect 46672 4320 46736 4324
rect 46752 4380 46816 4384
rect 46752 4324 46756 4380
rect 46756 4324 46812 4380
rect 46812 4324 46816 4380
rect 46752 4320 46816 4324
rect 46832 4380 46896 4384
rect 46832 4324 46836 4380
rect 46836 4324 46892 4380
rect 46892 4324 46896 4380
rect 46832 4320 46896 4324
rect 46912 4380 46976 4384
rect 46912 4324 46916 4380
rect 46916 4324 46972 4380
rect 46972 4324 46976 4380
rect 46912 4320 46976 4324
rect 6667 3836 6731 3840
rect 6667 3780 6671 3836
rect 6671 3780 6727 3836
rect 6727 3780 6731 3836
rect 6667 3776 6731 3780
rect 6747 3836 6811 3840
rect 6747 3780 6751 3836
rect 6751 3780 6807 3836
rect 6807 3780 6811 3836
rect 6747 3776 6811 3780
rect 6827 3836 6891 3840
rect 6827 3780 6831 3836
rect 6831 3780 6887 3836
rect 6887 3780 6891 3836
rect 6827 3776 6891 3780
rect 6907 3836 6971 3840
rect 6907 3780 6911 3836
rect 6911 3780 6967 3836
rect 6967 3780 6971 3836
rect 6907 3776 6971 3780
rect 18097 3836 18161 3840
rect 18097 3780 18101 3836
rect 18101 3780 18157 3836
rect 18157 3780 18161 3836
rect 18097 3776 18161 3780
rect 18177 3836 18241 3840
rect 18177 3780 18181 3836
rect 18181 3780 18237 3836
rect 18237 3780 18241 3836
rect 18177 3776 18241 3780
rect 18257 3836 18321 3840
rect 18257 3780 18261 3836
rect 18261 3780 18317 3836
rect 18317 3780 18321 3836
rect 18257 3776 18321 3780
rect 18337 3836 18401 3840
rect 18337 3780 18341 3836
rect 18341 3780 18397 3836
rect 18397 3780 18401 3836
rect 18337 3776 18401 3780
rect 29527 3836 29591 3840
rect 29527 3780 29531 3836
rect 29531 3780 29587 3836
rect 29587 3780 29591 3836
rect 29527 3776 29591 3780
rect 29607 3836 29671 3840
rect 29607 3780 29611 3836
rect 29611 3780 29667 3836
rect 29667 3780 29671 3836
rect 29607 3776 29671 3780
rect 29687 3836 29751 3840
rect 29687 3780 29691 3836
rect 29691 3780 29747 3836
rect 29747 3780 29751 3836
rect 29687 3776 29751 3780
rect 29767 3836 29831 3840
rect 29767 3780 29771 3836
rect 29771 3780 29827 3836
rect 29827 3780 29831 3836
rect 29767 3776 29831 3780
rect 40957 3836 41021 3840
rect 40957 3780 40961 3836
rect 40961 3780 41017 3836
rect 41017 3780 41021 3836
rect 40957 3776 41021 3780
rect 41037 3836 41101 3840
rect 41037 3780 41041 3836
rect 41041 3780 41097 3836
rect 41097 3780 41101 3836
rect 41037 3776 41101 3780
rect 41117 3836 41181 3840
rect 41117 3780 41121 3836
rect 41121 3780 41177 3836
rect 41177 3780 41181 3836
rect 41117 3776 41181 3780
rect 41197 3836 41261 3840
rect 41197 3780 41201 3836
rect 41201 3780 41257 3836
rect 41257 3780 41261 3836
rect 41197 3776 41261 3780
rect 12382 3292 12446 3296
rect 12382 3236 12386 3292
rect 12386 3236 12442 3292
rect 12442 3236 12446 3292
rect 12382 3232 12446 3236
rect 12462 3292 12526 3296
rect 12462 3236 12466 3292
rect 12466 3236 12522 3292
rect 12522 3236 12526 3292
rect 12462 3232 12526 3236
rect 12542 3292 12606 3296
rect 12542 3236 12546 3292
rect 12546 3236 12602 3292
rect 12602 3236 12606 3292
rect 12542 3232 12606 3236
rect 12622 3292 12686 3296
rect 12622 3236 12626 3292
rect 12626 3236 12682 3292
rect 12682 3236 12686 3292
rect 12622 3232 12686 3236
rect 23812 3292 23876 3296
rect 23812 3236 23816 3292
rect 23816 3236 23872 3292
rect 23872 3236 23876 3292
rect 23812 3232 23876 3236
rect 23892 3292 23956 3296
rect 23892 3236 23896 3292
rect 23896 3236 23952 3292
rect 23952 3236 23956 3292
rect 23892 3232 23956 3236
rect 23972 3292 24036 3296
rect 23972 3236 23976 3292
rect 23976 3236 24032 3292
rect 24032 3236 24036 3292
rect 23972 3232 24036 3236
rect 24052 3292 24116 3296
rect 24052 3236 24056 3292
rect 24056 3236 24112 3292
rect 24112 3236 24116 3292
rect 24052 3232 24116 3236
rect 35242 3292 35306 3296
rect 35242 3236 35246 3292
rect 35246 3236 35302 3292
rect 35302 3236 35306 3292
rect 35242 3232 35306 3236
rect 35322 3292 35386 3296
rect 35322 3236 35326 3292
rect 35326 3236 35382 3292
rect 35382 3236 35386 3292
rect 35322 3232 35386 3236
rect 35402 3292 35466 3296
rect 35402 3236 35406 3292
rect 35406 3236 35462 3292
rect 35462 3236 35466 3292
rect 35402 3232 35466 3236
rect 35482 3292 35546 3296
rect 35482 3236 35486 3292
rect 35486 3236 35542 3292
rect 35542 3236 35546 3292
rect 35482 3232 35546 3236
rect 46672 3292 46736 3296
rect 46672 3236 46676 3292
rect 46676 3236 46732 3292
rect 46732 3236 46736 3292
rect 46672 3232 46736 3236
rect 46752 3292 46816 3296
rect 46752 3236 46756 3292
rect 46756 3236 46812 3292
rect 46812 3236 46816 3292
rect 46752 3232 46816 3236
rect 46832 3292 46896 3296
rect 46832 3236 46836 3292
rect 46836 3236 46892 3292
rect 46892 3236 46896 3292
rect 46832 3232 46896 3236
rect 46912 3292 46976 3296
rect 46912 3236 46916 3292
rect 46916 3236 46972 3292
rect 46972 3236 46976 3292
rect 46912 3232 46976 3236
rect 6667 2748 6731 2752
rect 6667 2692 6671 2748
rect 6671 2692 6727 2748
rect 6727 2692 6731 2748
rect 6667 2688 6731 2692
rect 6747 2748 6811 2752
rect 6747 2692 6751 2748
rect 6751 2692 6807 2748
rect 6807 2692 6811 2748
rect 6747 2688 6811 2692
rect 6827 2748 6891 2752
rect 6827 2692 6831 2748
rect 6831 2692 6887 2748
rect 6887 2692 6891 2748
rect 6827 2688 6891 2692
rect 6907 2748 6971 2752
rect 6907 2692 6911 2748
rect 6911 2692 6967 2748
rect 6967 2692 6971 2748
rect 6907 2688 6971 2692
rect 18097 2748 18161 2752
rect 18097 2692 18101 2748
rect 18101 2692 18157 2748
rect 18157 2692 18161 2748
rect 18097 2688 18161 2692
rect 18177 2748 18241 2752
rect 18177 2692 18181 2748
rect 18181 2692 18237 2748
rect 18237 2692 18241 2748
rect 18177 2688 18241 2692
rect 18257 2748 18321 2752
rect 18257 2692 18261 2748
rect 18261 2692 18317 2748
rect 18317 2692 18321 2748
rect 18257 2688 18321 2692
rect 18337 2748 18401 2752
rect 18337 2692 18341 2748
rect 18341 2692 18397 2748
rect 18397 2692 18401 2748
rect 18337 2688 18401 2692
rect 29527 2748 29591 2752
rect 29527 2692 29531 2748
rect 29531 2692 29587 2748
rect 29587 2692 29591 2748
rect 29527 2688 29591 2692
rect 29607 2748 29671 2752
rect 29607 2692 29611 2748
rect 29611 2692 29667 2748
rect 29667 2692 29671 2748
rect 29607 2688 29671 2692
rect 29687 2748 29751 2752
rect 29687 2692 29691 2748
rect 29691 2692 29747 2748
rect 29747 2692 29751 2748
rect 29687 2688 29751 2692
rect 29767 2748 29831 2752
rect 29767 2692 29771 2748
rect 29771 2692 29827 2748
rect 29827 2692 29831 2748
rect 29767 2688 29831 2692
rect 40957 2748 41021 2752
rect 40957 2692 40961 2748
rect 40961 2692 41017 2748
rect 41017 2692 41021 2748
rect 40957 2688 41021 2692
rect 41037 2748 41101 2752
rect 41037 2692 41041 2748
rect 41041 2692 41097 2748
rect 41097 2692 41101 2748
rect 41037 2688 41101 2692
rect 41117 2748 41181 2752
rect 41117 2692 41121 2748
rect 41121 2692 41177 2748
rect 41177 2692 41181 2748
rect 41117 2688 41181 2692
rect 41197 2748 41261 2752
rect 41197 2692 41201 2748
rect 41201 2692 41257 2748
rect 41257 2692 41261 2748
rect 41197 2688 41261 2692
rect 12382 2204 12446 2208
rect 12382 2148 12386 2204
rect 12386 2148 12442 2204
rect 12442 2148 12446 2204
rect 12382 2144 12446 2148
rect 12462 2204 12526 2208
rect 12462 2148 12466 2204
rect 12466 2148 12522 2204
rect 12522 2148 12526 2204
rect 12462 2144 12526 2148
rect 12542 2204 12606 2208
rect 12542 2148 12546 2204
rect 12546 2148 12602 2204
rect 12602 2148 12606 2204
rect 12542 2144 12606 2148
rect 12622 2204 12686 2208
rect 12622 2148 12626 2204
rect 12626 2148 12682 2204
rect 12682 2148 12686 2204
rect 12622 2144 12686 2148
rect 23812 2204 23876 2208
rect 23812 2148 23816 2204
rect 23816 2148 23872 2204
rect 23872 2148 23876 2204
rect 23812 2144 23876 2148
rect 23892 2204 23956 2208
rect 23892 2148 23896 2204
rect 23896 2148 23952 2204
rect 23952 2148 23956 2204
rect 23892 2144 23956 2148
rect 23972 2204 24036 2208
rect 23972 2148 23976 2204
rect 23976 2148 24032 2204
rect 24032 2148 24036 2204
rect 23972 2144 24036 2148
rect 24052 2204 24116 2208
rect 24052 2148 24056 2204
rect 24056 2148 24112 2204
rect 24112 2148 24116 2204
rect 24052 2144 24116 2148
rect 35242 2204 35306 2208
rect 35242 2148 35246 2204
rect 35246 2148 35302 2204
rect 35302 2148 35306 2204
rect 35242 2144 35306 2148
rect 35322 2204 35386 2208
rect 35322 2148 35326 2204
rect 35326 2148 35382 2204
rect 35382 2148 35386 2204
rect 35322 2144 35386 2148
rect 35402 2204 35466 2208
rect 35402 2148 35406 2204
rect 35406 2148 35462 2204
rect 35462 2148 35466 2204
rect 35402 2144 35466 2148
rect 35482 2204 35546 2208
rect 35482 2148 35486 2204
rect 35486 2148 35542 2204
rect 35542 2148 35546 2204
rect 35482 2144 35546 2148
rect 46672 2204 46736 2208
rect 46672 2148 46676 2204
rect 46676 2148 46732 2204
rect 46732 2148 46736 2204
rect 46672 2144 46736 2148
rect 46752 2204 46816 2208
rect 46752 2148 46756 2204
rect 46756 2148 46812 2204
rect 46812 2148 46816 2204
rect 46752 2144 46816 2148
rect 46832 2204 46896 2208
rect 46832 2148 46836 2204
rect 46836 2148 46892 2204
rect 46892 2148 46896 2204
rect 46832 2144 46896 2148
rect 46912 2204 46976 2208
rect 46912 2148 46916 2204
rect 46916 2148 46972 2204
rect 46972 2148 46976 2204
rect 46912 2144 46976 2148
rect 6667 1660 6731 1664
rect 6667 1604 6671 1660
rect 6671 1604 6727 1660
rect 6727 1604 6731 1660
rect 6667 1600 6731 1604
rect 6747 1660 6811 1664
rect 6747 1604 6751 1660
rect 6751 1604 6807 1660
rect 6807 1604 6811 1660
rect 6747 1600 6811 1604
rect 6827 1660 6891 1664
rect 6827 1604 6831 1660
rect 6831 1604 6887 1660
rect 6887 1604 6891 1660
rect 6827 1600 6891 1604
rect 6907 1660 6971 1664
rect 6907 1604 6911 1660
rect 6911 1604 6967 1660
rect 6967 1604 6971 1660
rect 6907 1600 6971 1604
rect 18097 1660 18161 1664
rect 18097 1604 18101 1660
rect 18101 1604 18157 1660
rect 18157 1604 18161 1660
rect 18097 1600 18161 1604
rect 18177 1660 18241 1664
rect 18177 1604 18181 1660
rect 18181 1604 18237 1660
rect 18237 1604 18241 1660
rect 18177 1600 18241 1604
rect 18257 1660 18321 1664
rect 18257 1604 18261 1660
rect 18261 1604 18317 1660
rect 18317 1604 18321 1660
rect 18257 1600 18321 1604
rect 18337 1660 18401 1664
rect 18337 1604 18341 1660
rect 18341 1604 18397 1660
rect 18397 1604 18401 1660
rect 18337 1600 18401 1604
rect 29527 1660 29591 1664
rect 29527 1604 29531 1660
rect 29531 1604 29587 1660
rect 29587 1604 29591 1660
rect 29527 1600 29591 1604
rect 29607 1660 29671 1664
rect 29607 1604 29611 1660
rect 29611 1604 29667 1660
rect 29667 1604 29671 1660
rect 29607 1600 29671 1604
rect 29687 1660 29751 1664
rect 29687 1604 29691 1660
rect 29691 1604 29747 1660
rect 29747 1604 29751 1660
rect 29687 1600 29751 1604
rect 29767 1660 29831 1664
rect 29767 1604 29771 1660
rect 29771 1604 29827 1660
rect 29827 1604 29831 1660
rect 29767 1600 29831 1604
rect 40957 1660 41021 1664
rect 40957 1604 40961 1660
rect 40961 1604 41017 1660
rect 41017 1604 41021 1660
rect 40957 1600 41021 1604
rect 41037 1660 41101 1664
rect 41037 1604 41041 1660
rect 41041 1604 41097 1660
rect 41097 1604 41101 1660
rect 41037 1600 41101 1604
rect 41117 1660 41181 1664
rect 41117 1604 41121 1660
rect 41121 1604 41177 1660
rect 41177 1604 41181 1660
rect 41117 1600 41181 1604
rect 41197 1660 41261 1664
rect 41197 1604 41201 1660
rect 41201 1604 41257 1660
rect 41257 1604 41261 1660
rect 41197 1600 41261 1604
rect 12382 1116 12446 1120
rect 12382 1060 12386 1116
rect 12386 1060 12442 1116
rect 12442 1060 12446 1116
rect 12382 1056 12446 1060
rect 12462 1116 12526 1120
rect 12462 1060 12466 1116
rect 12466 1060 12522 1116
rect 12522 1060 12526 1116
rect 12462 1056 12526 1060
rect 12542 1116 12606 1120
rect 12542 1060 12546 1116
rect 12546 1060 12602 1116
rect 12602 1060 12606 1116
rect 12542 1056 12606 1060
rect 12622 1116 12686 1120
rect 12622 1060 12626 1116
rect 12626 1060 12682 1116
rect 12682 1060 12686 1116
rect 12622 1056 12686 1060
rect 23812 1116 23876 1120
rect 23812 1060 23816 1116
rect 23816 1060 23872 1116
rect 23872 1060 23876 1116
rect 23812 1056 23876 1060
rect 23892 1116 23956 1120
rect 23892 1060 23896 1116
rect 23896 1060 23952 1116
rect 23952 1060 23956 1116
rect 23892 1056 23956 1060
rect 23972 1116 24036 1120
rect 23972 1060 23976 1116
rect 23976 1060 24032 1116
rect 24032 1060 24036 1116
rect 23972 1056 24036 1060
rect 24052 1116 24116 1120
rect 24052 1060 24056 1116
rect 24056 1060 24112 1116
rect 24112 1060 24116 1116
rect 24052 1056 24116 1060
rect 35242 1116 35306 1120
rect 35242 1060 35246 1116
rect 35246 1060 35302 1116
rect 35302 1060 35306 1116
rect 35242 1056 35306 1060
rect 35322 1116 35386 1120
rect 35322 1060 35326 1116
rect 35326 1060 35382 1116
rect 35382 1060 35386 1116
rect 35322 1056 35386 1060
rect 35402 1116 35466 1120
rect 35402 1060 35406 1116
rect 35406 1060 35462 1116
rect 35462 1060 35466 1116
rect 35402 1056 35466 1060
rect 35482 1116 35546 1120
rect 35482 1060 35486 1116
rect 35486 1060 35542 1116
rect 35542 1060 35546 1116
rect 35482 1056 35546 1060
rect 46672 1116 46736 1120
rect 46672 1060 46676 1116
rect 46676 1060 46732 1116
rect 46732 1060 46736 1116
rect 46672 1056 46736 1060
rect 46752 1116 46816 1120
rect 46752 1060 46756 1116
rect 46756 1060 46812 1116
rect 46812 1060 46816 1116
rect 46752 1056 46816 1060
rect 46832 1116 46896 1120
rect 46832 1060 46836 1116
rect 46836 1060 46892 1116
rect 46892 1060 46896 1116
rect 46832 1056 46896 1060
rect 46912 1116 46976 1120
rect 46912 1060 46916 1116
rect 46916 1060 46972 1116
rect 46972 1060 46976 1116
rect 46912 1056 46976 1060
<< metal4 >>
rect 6659 8192 6979 8752
rect 6659 8128 6667 8192
rect 6731 8128 6747 8192
rect 6811 8128 6827 8192
rect 6891 8128 6907 8192
rect 6971 8128 6979 8192
rect 6659 7104 6979 8128
rect 6659 7040 6667 7104
rect 6731 7040 6747 7104
rect 6811 7040 6827 7104
rect 6891 7040 6907 7104
rect 6971 7040 6979 7104
rect 6659 6016 6979 7040
rect 6659 5952 6667 6016
rect 6731 5952 6747 6016
rect 6811 5952 6827 6016
rect 6891 5952 6907 6016
rect 6971 5952 6979 6016
rect 6659 4928 6979 5952
rect 6659 4864 6667 4928
rect 6731 4864 6747 4928
rect 6811 4864 6827 4928
rect 6891 4864 6907 4928
rect 6971 4864 6979 4928
rect 6659 3840 6979 4864
rect 6659 3776 6667 3840
rect 6731 3776 6747 3840
rect 6811 3776 6827 3840
rect 6891 3776 6907 3840
rect 6971 3776 6979 3840
rect 6659 2752 6979 3776
rect 6659 2688 6667 2752
rect 6731 2688 6747 2752
rect 6811 2688 6827 2752
rect 6891 2688 6907 2752
rect 6971 2688 6979 2752
rect 6659 1664 6979 2688
rect 6659 1600 6667 1664
rect 6731 1600 6747 1664
rect 6811 1600 6827 1664
rect 6891 1600 6907 1664
rect 6971 1600 6979 1664
rect 6659 1040 6979 1600
rect 12374 8736 12694 8752
rect 12374 8672 12382 8736
rect 12446 8672 12462 8736
rect 12526 8672 12542 8736
rect 12606 8672 12622 8736
rect 12686 8672 12694 8736
rect 12374 7648 12694 8672
rect 12374 7584 12382 7648
rect 12446 7584 12462 7648
rect 12526 7584 12542 7648
rect 12606 7584 12622 7648
rect 12686 7584 12694 7648
rect 12374 6560 12694 7584
rect 12374 6496 12382 6560
rect 12446 6496 12462 6560
rect 12526 6496 12542 6560
rect 12606 6496 12622 6560
rect 12686 6496 12694 6560
rect 12374 5472 12694 6496
rect 12374 5408 12382 5472
rect 12446 5408 12462 5472
rect 12526 5408 12542 5472
rect 12606 5408 12622 5472
rect 12686 5408 12694 5472
rect 12374 4384 12694 5408
rect 12374 4320 12382 4384
rect 12446 4320 12462 4384
rect 12526 4320 12542 4384
rect 12606 4320 12622 4384
rect 12686 4320 12694 4384
rect 12374 3296 12694 4320
rect 12374 3232 12382 3296
rect 12446 3232 12462 3296
rect 12526 3232 12542 3296
rect 12606 3232 12622 3296
rect 12686 3232 12694 3296
rect 12374 2208 12694 3232
rect 12374 2144 12382 2208
rect 12446 2144 12462 2208
rect 12526 2144 12542 2208
rect 12606 2144 12622 2208
rect 12686 2144 12694 2208
rect 12374 1120 12694 2144
rect 12374 1056 12382 1120
rect 12446 1056 12462 1120
rect 12526 1056 12542 1120
rect 12606 1056 12622 1120
rect 12686 1056 12694 1120
rect 12374 1040 12694 1056
rect 18089 8192 18409 8752
rect 18089 8128 18097 8192
rect 18161 8128 18177 8192
rect 18241 8128 18257 8192
rect 18321 8128 18337 8192
rect 18401 8128 18409 8192
rect 18089 7104 18409 8128
rect 18089 7040 18097 7104
rect 18161 7040 18177 7104
rect 18241 7040 18257 7104
rect 18321 7040 18337 7104
rect 18401 7040 18409 7104
rect 18089 6016 18409 7040
rect 18089 5952 18097 6016
rect 18161 5952 18177 6016
rect 18241 5952 18257 6016
rect 18321 5952 18337 6016
rect 18401 5952 18409 6016
rect 18089 4928 18409 5952
rect 18089 4864 18097 4928
rect 18161 4864 18177 4928
rect 18241 4864 18257 4928
rect 18321 4864 18337 4928
rect 18401 4864 18409 4928
rect 18089 3840 18409 4864
rect 18089 3776 18097 3840
rect 18161 3776 18177 3840
rect 18241 3776 18257 3840
rect 18321 3776 18337 3840
rect 18401 3776 18409 3840
rect 18089 2752 18409 3776
rect 18089 2688 18097 2752
rect 18161 2688 18177 2752
rect 18241 2688 18257 2752
rect 18321 2688 18337 2752
rect 18401 2688 18409 2752
rect 18089 1664 18409 2688
rect 18089 1600 18097 1664
rect 18161 1600 18177 1664
rect 18241 1600 18257 1664
rect 18321 1600 18337 1664
rect 18401 1600 18409 1664
rect 18089 1040 18409 1600
rect 23804 8736 24124 8752
rect 23804 8672 23812 8736
rect 23876 8672 23892 8736
rect 23956 8672 23972 8736
rect 24036 8672 24052 8736
rect 24116 8672 24124 8736
rect 23804 7648 24124 8672
rect 23804 7584 23812 7648
rect 23876 7584 23892 7648
rect 23956 7584 23972 7648
rect 24036 7584 24052 7648
rect 24116 7584 24124 7648
rect 23804 6560 24124 7584
rect 23804 6496 23812 6560
rect 23876 6496 23892 6560
rect 23956 6496 23972 6560
rect 24036 6496 24052 6560
rect 24116 6496 24124 6560
rect 23804 5472 24124 6496
rect 23804 5408 23812 5472
rect 23876 5408 23892 5472
rect 23956 5408 23972 5472
rect 24036 5408 24052 5472
rect 24116 5408 24124 5472
rect 23804 4384 24124 5408
rect 23804 4320 23812 4384
rect 23876 4320 23892 4384
rect 23956 4320 23972 4384
rect 24036 4320 24052 4384
rect 24116 4320 24124 4384
rect 23804 3296 24124 4320
rect 23804 3232 23812 3296
rect 23876 3232 23892 3296
rect 23956 3232 23972 3296
rect 24036 3232 24052 3296
rect 24116 3232 24124 3296
rect 23804 2208 24124 3232
rect 23804 2144 23812 2208
rect 23876 2144 23892 2208
rect 23956 2144 23972 2208
rect 24036 2144 24052 2208
rect 24116 2144 24124 2208
rect 23804 1120 24124 2144
rect 23804 1056 23812 1120
rect 23876 1056 23892 1120
rect 23956 1056 23972 1120
rect 24036 1056 24052 1120
rect 24116 1056 24124 1120
rect 23804 1040 24124 1056
rect 29519 8192 29839 8752
rect 29519 8128 29527 8192
rect 29591 8128 29607 8192
rect 29671 8128 29687 8192
rect 29751 8128 29767 8192
rect 29831 8128 29839 8192
rect 29519 7104 29839 8128
rect 29519 7040 29527 7104
rect 29591 7040 29607 7104
rect 29671 7040 29687 7104
rect 29751 7040 29767 7104
rect 29831 7040 29839 7104
rect 29519 6016 29839 7040
rect 29519 5952 29527 6016
rect 29591 5952 29607 6016
rect 29671 5952 29687 6016
rect 29751 5952 29767 6016
rect 29831 5952 29839 6016
rect 29519 4928 29839 5952
rect 29519 4864 29527 4928
rect 29591 4864 29607 4928
rect 29671 4864 29687 4928
rect 29751 4864 29767 4928
rect 29831 4864 29839 4928
rect 29519 3840 29839 4864
rect 29519 3776 29527 3840
rect 29591 3776 29607 3840
rect 29671 3776 29687 3840
rect 29751 3776 29767 3840
rect 29831 3776 29839 3840
rect 29519 2752 29839 3776
rect 29519 2688 29527 2752
rect 29591 2688 29607 2752
rect 29671 2688 29687 2752
rect 29751 2688 29767 2752
rect 29831 2688 29839 2752
rect 29519 1664 29839 2688
rect 29519 1600 29527 1664
rect 29591 1600 29607 1664
rect 29671 1600 29687 1664
rect 29751 1600 29767 1664
rect 29831 1600 29839 1664
rect 29519 1040 29839 1600
rect 35234 8736 35554 8752
rect 35234 8672 35242 8736
rect 35306 8672 35322 8736
rect 35386 8672 35402 8736
rect 35466 8672 35482 8736
rect 35546 8672 35554 8736
rect 35234 7648 35554 8672
rect 35234 7584 35242 7648
rect 35306 7584 35322 7648
rect 35386 7584 35402 7648
rect 35466 7584 35482 7648
rect 35546 7584 35554 7648
rect 35234 6560 35554 7584
rect 35234 6496 35242 6560
rect 35306 6496 35322 6560
rect 35386 6496 35402 6560
rect 35466 6496 35482 6560
rect 35546 6496 35554 6560
rect 35234 5472 35554 6496
rect 35234 5408 35242 5472
rect 35306 5408 35322 5472
rect 35386 5408 35402 5472
rect 35466 5408 35482 5472
rect 35546 5408 35554 5472
rect 35234 4384 35554 5408
rect 35234 4320 35242 4384
rect 35306 4320 35322 4384
rect 35386 4320 35402 4384
rect 35466 4320 35482 4384
rect 35546 4320 35554 4384
rect 35234 3296 35554 4320
rect 35234 3232 35242 3296
rect 35306 3232 35322 3296
rect 35386 3232 35402 3296
rect 35466 3232 35482 3296
rect 35546 3232 35554 3296
rect 35234 2208 35554 3232
rect 35234 2144 35242 2208
rect 35306 2144 35322 2208
rect 35386 2144 35402 2208
rect 35466 2144 35482 2208
rect 35546 2144 35554 2208
rect 35234 1120 35554 2144
rect 35234 1056 35242 1120
rect 35306 1056 35322 1120
rect 35386 1056 35402 1120
rect 35466 1056 35482 1120
rect 35546 1056 35554 1120
rect 35234 1040 35554 1056
rect 40949 8192 41269 8752
rect 40949 8128 40957 8192
rect 41021 8128 41037 8192
rect 41101 8128 41117 8192
rect 41181 8128 41197 8192
rect 41261 8128 41269 8192
rect 40949 7104 41269 8128
rect 40949 7040 40957 7104
rect 41021 7040 41037 7104
rect 41101 7040 41117 7104
rect 41181 7040 41197 7104
rect 41261 7040 41269 7104
rect 40949 6016 41269 7040
rect 40949 5952 40957 6016
rect 41021 5952 41037 6016
rect 41101 5952 41117 6016
rect 41181 5952 41197 6016
rect 41261 5952 41269 6016
rect 40949 4928 41269 5952
rect 40949 4864 40957 4928
rect 41021 4864 41037 4928
rect 41101 4864 41117 4928
rect 41181 4864 41197 4928
rect 41261 4864 41269 4928
rect 40949 3840 41269 4864
rect 40949 3776 40957 3840
rect 41021 3776 41037 3840
rect 41101 3776 41117 3840
rect 41181 3776 41197 3840
rect 41261 3776 41269 3840
rect 40949 2752 41269 3776
rect 40949 2688 40957 2752
rect 41021 2688 41037 2752
rect 41101 2688 41117 2752
rect 41181 2688 41197 2752
rect 41261 2688 41269 2752
rect 40949 1664 41269 2688
rect 40949 1600 40957 1664
rect 41021 1600 41037 1664
rect 41101 1600 41117 1664
rect 41181 1600 41197 1664
rect 41261 1600 41269 1664
rect 40949 1040 41269 1600
rect 46664 8736 46984 8752
rect 46664 8672 46672 8736
rect 46736 8672 46752 8736
rect 46816 8672 46832 8736
rect 46896 8672 46912 8736
rect 46976 8672 46984 8736
rect 46664 7648 46984 8672
rect 46664 7584 46672 7648
rect 46736 7584 46752 7648
rect 46816 7584 46832 7648
rect 46896 7584 46912 7648
rect 46976 7584 46984 7648
rect 46664 6560 46984 7584
rect 46664 6496 46672 6560
rect 46736 6496 46752 6560
rect 46816 6496 46832 6560
rect 46896 6496 46912 6560
rect 46976 6496 46984 6560
rect 46664 5472 46984 6496
rect 46664 5408 46672 5472
rect 46736 5408 46752 5472
rect 46816 5408 46832 5472
rect 46896 5408 46912 5472
rect 46976 5408 46984 5472
rect 46664 4384 46984 5408
rect 46664 4320 46672 4384
rect 46736 4320 46752 4384
rect 46816 4320 46832 4384
rect 46896 4320 46912 4384
rect 46976 4320 46984 4384
rect 46664 3296 46984 4320
rect 46664 3232 46672 3296
rect 46736 3232 46752 3296
rect 46816 3232 46832 3296
rect 46896 3232 46912 3296
rect 46976 3232 46984 3296
rect 46664 2208 46984 3232
rect 46664 2144 46672 2208
rect 46736 2144 46752 2208
rect 46816 2144 46832 2208
rect 46896 2144 46912 2208
rect 46976 2144 46984 2208
rect 46664 1120 46984 2144
rect 46664 1056 46672 1120
rect 46736 1056 46752 1120
rect 46816 1056 46832 1120
rect 46896 1056 46912 1120
rect 46976 1056 46984 1120
rect 46664 1040 46984 1056
use sky130_fd_sc_hd__decap_6  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_36
timestamp 1688980957
transform 1 0 4416 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_60
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_72
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_80 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_108
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_132
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_156
timestamp 1688980957
transform 1 0 15456 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_180
timestamp 1688980957
transform 1 0 17664 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_192
timestamp 1688980957
transform 1 0 18768 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_204
timestamp 1688980957
transform 1 0 19872 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_216
timestamp 1688980957
transform 1 0 20976 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_228
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_246 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_276
timestamp 1688980957
transform 1 0 26496 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_300
timestamp 1688980957
transform 1 0 28704 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_324
timestamp 1688980957
transform 1 0 30912 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_348
timestamp 1688980957
transform 1 0 33120 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_360
timestamp 1688980957
transform 1 0 34224 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_372
timestamp 1688980957
transform 1 0 35328 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_384
timestamp 1688980957
transform 1 0 36432 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_396
timestamp 1688980957
transform 1 0 37536 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_408
timestamp 1688980957
transform 1 0 38640 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_416
timestamp 1688980957
transform 1 0 39376 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_444
timestamp 1688980957
transform 1 0 41952 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_468
timestamp 1688980957
transform 1 0 44160 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_477
timestamp 1688980957
transform 1 0 44988 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_492 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46368 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_209
timestamp 1688980957
transform 1 0 20332 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_221
timestamp 1688980957
transform 1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_235
timestamp 1688980957
transform 1 0 22724 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_252
timestamp 1688980957
transform 1 0 24288 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_260
timestamp 1688980957
transform 1 0 25024 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_272
timestamp 1688980957
transform 1 0 26128 0 -1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_284
timestamp 1688980957
transform 1 0 27232 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_296
timestamp 1688980957
transform 1 0 28336 0 -1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_307
timestamp 1688980957
transform 1 0 29348 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_319
timestamp 1688980957
transform 1 0 30452 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_330
timestamp 1688980957
transform 1 0 31464 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_355
timestamp 1688980957
transform 1 0 33764 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_367
timestamp 1688980957
transform 1 0 34868 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_377
timestamp 1688980957
transform 1 0 35788 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_389
timestamp 1688980957
transform 1 0 36892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_397
timestamp 1688980957
transform 1 0 37628 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_401
timestamp 1688980957
transform 1 0 37996 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_413
timestamp 1688980957
transform 1 0 39100 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_425
timestamp 1688980957
transform 1 0 40204 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_437
timestamp 1688980957
transform 1 0 41308 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_445
timestamp 1688980957
transform 1 0 42044 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_452
timestamp 1688980957
transform 1 0 42688 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_464
timestamp 1688980957
transform 1 0 43792 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_470
timestamp 1688980957
transform 1 0 44344 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_475
timestamp 1688980957
transform 1 0 44804 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_483
timestamp 1688980957
transform 1 0 45540 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_487
timestamp 1688980957
transform 1 0 45908 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_493
timestamp 1688980957
transform 1 0 46460 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_220
timestamp 1688980957
transform 1 0 21344 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_232
timestamp 1688980957
transform 1 0 22448 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_238
timestamp 1688980957
transform 1 0 23000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_267
timestamp 1688980957
transform 1 0 25668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_290
timestamp 1688980957
transform 1 0 27784 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_302
timestamp 1688980957
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_314
timestamp 1688980957
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_326
timestamp 1688980957
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_334
timestamp 1688980957
transform 1 0 31832 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_338
timestamp 1688980957
transform 1 0 32200 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_350
timestamp 1688980957
transform 1 0 33304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_358
timestamp 1688980957
transform 1 0 34040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_362
timestamp 1688980957
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_383
timestamp 1688980957
transform 1 0 36340 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_387
timestamp 1688980957
transform 1 0 36708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_399
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_407
timestamp 1688980957
transform 1 0 38548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_411
timestamp 1688980957
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_453
timestamp 1688980957
transform 1 0 42780 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_459
timestamp 1688980957
transform 1 0 43332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_471
timestamp 1688980957
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1688980957
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_480
timestamp 1688980957
transform 1 0 45264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_488
timestamp 1688980957
transform 1 0 46000 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_485
timestamp 1688980957
transform 1 0 45724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_493
timestamp 1688980957
transform 1 0 46460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_489
timestamp 1688980957
transform 1 0 46092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_493
timestamp 1688980957
transform 1 0 46460 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_485
timestamp 1688980957
transform 1 0 45724 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_493
timestamp 1688980957
transform 1 0 46460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_489
timestamp 1688980957
transform 1 0 46092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_493
timestamp 1688980957
transform 1 0 46460 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_485
timestamp 1688980957
transform 1 0 45724 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_493
timestamp 1688980957
transform 1 0 46460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_489
timestamp 1688980957
transform 1 0 46092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_493
timestamp 1688980957
transform 1 0 46460 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_485
timestamp 1688980957
transform 1 0 45724 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_493
timestamp 1688980957
transform 1 0 46460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_481
timestamp 1688980957
transform 1 0 45356 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_21
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_33
timestamp 1688980957
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_204
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_208
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_215
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_236
timestamp 1688980957
transform 1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_248
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_252
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_259
timestamp 1688980957
transform 1 0 24932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_271
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_469
timestamp 1688980957
transform 1 0 44252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_17
timestamp 1688980957
transform 1 0 2668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1688980957
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_69
timestamp 1688980957
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1688980957
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_100
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_112
timestamp 1688980957
transform 1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_128
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_160
timestamp 1688980957
transform 1 0 15824 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_176
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_180
timestamp 1688980957
transform 1 0 17664 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_260
timestamp 1688980957
transform 1 0 25024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_288
timestamp 1688980957
transform 1 0 27600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_292
timestamp 1688980957
transform 1 0 27968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_296
timestamp 1688980957
transform 1 0 28336 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_300
timestamp 1688980957
transform 1 0 28704 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_304
timestamp 1688980957
transform 1 0 29072 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_313
timestamp 1688980957
transform 1 0 29900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_325
timestamp 1688980957
transform 1 0 31004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_337
timestamp 1688980957
transform 1 0 32108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_349
timestamp 1688980957
transform 1 0 33212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_361
timestamp 1688980957
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_437
timestamp 1688980957
transform 1 0 41308 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_449
timestamp 1688980957
transform 1 0 42412 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_463
timestamp 1688980957
transform 1 0 43700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_471
timestamp 1688980957
transform 1 0 44436 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_489
timestamp 1688980957
transform 1 0 46092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_493
timestamp 1688980957
transform 1 0 46460 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_89
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_124
timestamp 1688980957
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_156
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_203
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_213
timestamp 1688980957
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_256
timestamp 1688980957
transform 1 0 24656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_260
timestamp 1688980957
transform 1 0 25024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_264
timestamp 1688980957
transform 1 0 25392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_268
timestamp 1688980957
transform 1 0 25760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_272
timestamp 1688980957
transform 1 0 26128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_276
timestamp 1688980957
transform 1 0 26496 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_284
timestamp 1688980957
transform 1 0 27232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_288
timestamp 1688980957
transform 1 0 27600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_292
timestamp 1688980957
transform 1 0 27968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_296
timestamp 1688980957
transform 1 0 28336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_300
timestamp 1688980957
transform 1 0 28704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_304
timestamp 1688980957
transform 1 0 29072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_312
timestamp 1688980957
transform 1 0 29808 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_316
timestamp 1688980957
transform 1 0 30176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_320
timestamp 1688980957
transform 1 0 30544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_324
timestamp 1688980957
transform 1 0 30912 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_328
timestamp 1688980957
transform 1 0 31280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_332
timestamp 1688980957
transform 1 0 31648 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_340
timestamp 1688980957
transform 1 0 32384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_344
timestamp 1688980957
transform 1 0 32752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_348
timestamp 1688980957
transform 1 0 33120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_352
timestamp 1688980957
transform 1 0 33488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_356
timestamp 1688980957
transform 1 0 33856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_360
timestamp 1688980957
transform 1 0 34224 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_368
timestamp 1688980957
transform 1 0 34960 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_372
timestamp 1688980957
transform 1 0 35328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_376
timestamp 1688980957
transform 1 0 35696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_380
timestamp 1688980957
transform 1 0 36064 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_384
timestamp 1688980957
transform 1 0 36432 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_388
timestamp 1688980957
transform 1 0 36800 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_396
timestamp 1688980957
transform 1 0 37536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_400
timestamp 1688980957
transform 1 0 37904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_404
timestamp 1688980957
transform 1 0 38272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_408
timestamp 1688980957
transform 1 0 38640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_412
timestamp 1688980957
transform 1 0 39008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_416
timestamp 1688980957
transform 1 0 39376 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_443
timestamp 1688980957
transform 1 0 41860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_473
timestamp 1688980957
transform 1 0 44620 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_489
timestamp 1688980957
transform 1 0 46092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_493
timestamp 1688980957
transform 1 0 46460 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26496 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 28704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 30912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 33120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 35328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 37536 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 39744 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 41952 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 44160 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 46092 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 10764 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 12972 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform -1 0 15456 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform -1 0 17664 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 19872 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform -1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform -1 0 24288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 19596 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform -1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 24748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 27324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 27692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform -1 0 32016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform -1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 32476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform -1 0 33120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform -1 0 33488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 28428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 28796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 29900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 30636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 31004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform -1 0 33856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform -1 0 37536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform -1 0 37904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform -1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform -1 0 38640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform -1 0 39008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform -1 0 39376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform -1 0 34224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1688980957
transform -1 0 34592 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform -1 0 34960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform -1 0 35328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform -1 0 35696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1688980957
transform -1 0 36064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform -1 0 36432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1688980957
transform -1 0 36800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1688980957
transform -1 0 37168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform 1 0 1932 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  inst_clk_buf
timestamp 1688980957
transform 1 0 24748 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__00_
timestamp 1688980957
transform -1 0 27048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__01_
timestamp 1688980957
transform -1 0 26772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__02_
timestamp 1688980957
transform -1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__03_
timestamp 1688980957
transform -1 0 26220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__04_
timestamp 1688980957
transform -1 0 25392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__05_
timestamp 1688980957
transform -1 0 25024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__06_
timestamp 1688980957
transform -1 0 24288 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__07_
timestamp 1688980957
transform -1 0 24288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__08_
timestamp 1688980957
transform -1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__09_
timestamp 1688980957
transform -1 0 22632 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__10_
timestamp 1688980957
transform -1 0 22356 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__11_
timestamp 1688980957
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__12_
timestamp 1688980957
transform -1 0 22080 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__13_
timestamp 1688980957
transform -1 0 21804 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__14_
timestamp 1688980957
transform -1 0 21528 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__15_
timestamp 1688980957
transform -1 0 21252 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__16_
timestamp 1688980957
transform -1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__17_
timestamp 1688980957
transform -1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__18_
timestamp 1688980957
transform -1 0 29072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__19_
timestamp 1688980957
transform -1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__20_
timestamp 1688980957
transform -1 0 28336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__21_
timestamp 1688980957
transform -1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__22_
timestamp 1688980957
transform -1 0 27600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__23_
timestamp 1688980957
transform -1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__24_
timestamp 1688980957
transform -1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__25_
timestamp 1688980957
transform -1 0 24656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__26_
timestamp 1688980957
transform -1 0 24748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__27_
timestamp 1688980957
transform -1 0 24932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__28_
timestamp 1688980957
transform -1 0 25944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__29_
timestamp 1688980957
transform -1 0 25668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__30_
timestamp 1688980957
transform -1 0 29900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__31_
timestamp 1688980957
transform -1 0 29440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__32_
timestamp 1688980957
transform -1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__33_
timestamp 1688980957
transform 1 0 22632 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__34_
timestamp 1688980957
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__35_
timestamp 1688980957
transform 1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__36_
timestamp 1688980957
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__37_
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__38_
timestamp 1688980957
transform -1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__39_
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__40_
timestamp 1688980957
transform -1 0 23736 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__41_
timestamp 1688980957
transform 1 0 22908 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__42_
timestamp 1688980957
transform 1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__43_
timestamp 1688980957
transform 1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__44_
timestamp 1688980957
transform 1 0 23092 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__45_
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__46_
timestamp 1688980957
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__47_
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__48_
timestamp 1688980957
transform -1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__49_
timestamp 1688980957
transform -1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__50_
timestamp 1688980957
transform -1 0 19596 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__51_
timestamp 1688980957
transform -1 0 19136 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 43884 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 45540 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 44896 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 45448 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 44344 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 45448 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 46000 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 46000 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 45540 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 41308 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 42964 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 44068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 44988 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform -1 0 2300 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform -1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform -1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1688980957
transform -1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform -1 0 2944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1688980957
transform -1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform -1 0 4508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform -1 0 4416 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1688980957
transform -1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1688980957
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform -1 0 5336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform -1 0 5888 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform -1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform -1 0 6992 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1688980957
transform -1 0 7452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1688980957
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform -1 0 8280 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1688980957
transform -1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform -1 0 12512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1688980957
transform -1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1688980957
transform -1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1688980957
transform -1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform -1 0 13984 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1688980957
transform -1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform -1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform -1 0 8832 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform -1 0 9936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1688980957
transform -1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1688980957
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform -1 0 11408 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform -1 0 12236 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 17848 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1688980957
transform 1 0 18400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1688980957
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform -1 0 19780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1688980957
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1688980957
transform -1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform -1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform -1 0 15456 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1688980957
transform -1 0 15824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1688980957
transform -1 0 16008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform -1 0 16560 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1688980957
transform -1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1688980957
transform -1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform -1 0 17848 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 46828 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 46828 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 46828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 46828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 46828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 46828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 46828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 46828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 46828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 46828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 46828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 46828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 46828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform -1 0 23736 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform -1 0 23184 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform -1 0 23460 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform -1 0 24012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform -1 0 23736 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform -1 0 23460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform -1 0 22448 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform -1 0 20332 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform -1 0 22724 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform -1 0 24748 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform -1 0 27232 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform -1 0 29348 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform -1 0 31464 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform -1 0 33764 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform -1 0 35788 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform -1 0 37996 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform -1 0 44344 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform -1 0 42688 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform -1 0 44804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform -1 0 45908 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 25116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 24012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_7__0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 23092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 25392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 31924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 34132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 38640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform -1 0 45724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 45724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 44896 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 4066 0 4122 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 26146 0 26202 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 28354 0 28410 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 30562 0 30618 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 32770 0 32826 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 34978 0 35034 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 37186 0 37242 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 39394 0 39450 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 41602 0 41658 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 43810 0 43866 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 46018 0 46074 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 39762 9840 39818 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 43442 9840 43498 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 43810 9840 43866 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 44178 9840 44234 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 44546 9840 44602 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 44914 9840 44970 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 45282 9840 45338 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 45650 9840 45706 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 46018 9840 46074 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 46386 9840 46442 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 46754 9840 46810 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 40130 9840 40186 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 40498 9840 40554 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 40866 9840 40922 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 41234 9840 41290 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 41602 9840 41658 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 41970 9840 42026 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 42338 9840 42394 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 42706 9840 42762 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 43074 9840 43130 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 1122 9840 1178 10000 0 FreeSans 224 90 0 0 N1BEG[0]
port 40 nsew signal tristate
flabel metal2 s 1490 9840 1546 10000 0 FreeSans 224 90 0 0 N1BEG[1]
port 41 nsew signal tristate
flabel metal2 s 1858 9840 1914 10000 0 FreeSans 224 90 0 0 N1BEG[2]
port 42 nsew signal tristate
flabel metal2 s 2226 9840 2282 10000 0 FreeSans 224 90 0 0 N1BEG[3]
port 43 nsew signal tristate
flabel metal2 s 2594 9840 2650 10000 0 FreeSans 224 90 0 0 N2BEG[0]
port 44 nsew signal tristate
flabel metal2 s 2962 9840 3018 10000 0 FreeSans 224 90 0 0 N2BEG[1]
port 45 nsew signal tristate
flabel metal2 s 3330 9840 3386 10000 0 FreeSans 224 90 0 0 N2BEG[2]
port 46 nsew signal tristate
flabel metal2 s 3698 9840 3754 10000 0 FreeSans 224 90 0 0 N2BEG[3]
port 47 nsew signal tristate
flabel metal2 s 4066 9840 4122 10000 0 FreeSans 224 90 0 0 N2BEG[4]
port 48 nsew signal tristate
flabel metal2 s 4434 9840 4490 10000 0 FreeSans 224 90 0 0 N2BEG[5]
port 49 nsew signal tristate
flabel metal2 s 4802 9840 4858 10000 0 FreeSans 224 90 0 0 N2BEG[6]
port 50 nsew signal tristate
flabel metal2 s 5170 9840 5226 10000 0 FreeSans 224 90 0 0 N2BEG[7]
port 51 nsew signal tristate
flabel metal2 s 5538 9840 5594 10000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 52 nsew signal tristate
flabel metal2 s 5906 9840 5962 10000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 53 nsew signal tristate
flabel metal2 s 6274 9840 6330 10000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 54 nsew signal tristate
flabel metal2 s 6642 9840 6698 10000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 55 nsew signal tristate
flabel metal2 s 7010 9840 7066 10000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 56 nsew signal tristate
flabel metal2 s 7378 9840 7434 10000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 57 nsew signal tristate
flabel metal2 s 7746 9840 7802 10000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 58 nsew signal tristate
flabel metal2 s 8114 9840 8170 10000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 59 nsew signal tristate
flabel metal2 s 8482 9840 8538 10000 0 FreeSans 224 90 0 0 N4BEG[0]
port 60 nsew signal tristate
flabel metal2 s 12162 9840 12218 10000 0 FreeSans 224 90 0 0 N4BEG[10]
port 61 nsew signal tristate
flabel metal2 s 12530 9840 12586 10000 0 FreeSans 224 90 0 0 N4BEG[11]
port 62 nsew signal tristate
flabel metal2 s 12898 9840 12954 10000 0 FreeSans 224 90 0 0 N4BEG[12]
port 63 nsew signal tristate
flabel metal2 s 13266 9840 13322 10000 0 FreeSans 224 90 0 0 N4BEG[13]
port 64 nsew signal tristate
flabel metal2 s 13634 9840 13690 10000 0 FreeSans 224 90 0 0 N4BEG[14]
port 65 nsew signal tristate
flabel metal2 s 14002 9840 14058 10000 0 FreeSans 224 90 0 0 N4BEG[15]
port 66 nsew signal tristate
flabel metal2 s 8850 9840 8906 10000 0 FreeSans 224 90 0 0 N4BEG[1]
port 67 nsew signal tristate
flabel metal2 s 9218 9840 9274 10000 0 FreeSans 224 90 0 0 N4BEG[2]
port 68 nsew signal tristate
flabel metal2 s 9586 9840 9642 10000 0 FreeSans 224 90 0 0 N4BEG[3]
port 69 nsew signal tristate
flabel metal2 s 9954 9840 10010 10000 0 FreeSans 224 90 0 0 N4BEG[4]
port 70 nsew signal tristate
flabel metal2 s 10322 9840 10378 10000 0 FreeSans 224 90 0 0 N4BEG[5]
port 71 nsew signal tristate
flabel metal2 s 10690 9840 10746 10000 0 FreeSans 224 90 0 0 N4BEG[6]
port 72 nsew signal tristate
flabel metal2 s 11058 9840 11114 10000 0 FreeSans 224 90 0 0 N4BEG[7]
port 73 nsew signal tristate
flabel metal2 s 11426 9840 11482 10000 0 FreeSans 224 90 0 0 N4BEG[8]
port 74 nsew signal tristate
flabel metal2 s 11794 9840 11850 10000 0 FreeSans 224 90 0 0 N4BEG[9]
port 75 nsew signal tristate
flabel metal2 s 14370 9840 14426 10000 0 FreeSans 224 90 0 0 NN4BEG[0]
port 76 nsew signal tristate
flabel metal2 s 18050 9840 18106 10000 0 FreeSans 224 90 0 0 NN4BEG[10]
port 77 nsew signal tristate
flabel metal2 s 18418 9840 18474 10000 0 FreeSans 224 90 0 0 NN4BEG[11]
port 78 nsew signal tristate
flabel metal2 s 18786 9840 18842 10000 0 FreeSans 224 90 0 0 NN4BEG[12]
port 79 nsew signal tristate
flabel metal2 s 19154 9840 19210 10000 0 FreeSans 224 90 0 0 NN4BEG[13]
port 80 nsew signal tristate
flabel metal2 s 19522 9840 19578 10000 0 FreeSans 224 90 0 0 NN4BEG[14]
port 81 nsew signal tristate
flabel metal2 s 19890 9840 19946 10000 0 FreeSans 224 90 0 0 NN4BEG[15]
port 82 nsew signal tristate
flabel metal2 s 14738 9840 14794 10000 0 FreeSans 224 90 0 0 NN4BEG[1]
port 83 nsew signal tristate
flabel metal2 s 15106 9840 15162 10000 0 FreeSans 224 90 0 0 NN4BEG[2]
port 84 nsew signal tristate
flabel metal2 s 15474 9840 15530 10000 0 FreeSans 224 90 0 0 NN4BEG[3]
port 85 nsew signal tristate
flabel metal2 s 15842 9840 15898 10000 0 FreeSans 224 90 0 0 NN4BEG[4]
port 86 nsew signal tristate
flabel metal2 s 16210 9840 16266 10000 0 FreeSans 224 90 0 0 NN4BEG[5]
port 87 nsew signal tristate
flabel metal2 s 16578 9840 16634 10000 0 FreeSans 224 90 0 0 NN4BEG[6]
port 88 nsew signal tristate
flabel metal2 s 16946 9840 17002 10000 0 FreeSans 224 90 0 0 NN4BEG[7]
port 89 nsew signal tristate
flabel metal2 s 17314 9840 17370 10000 0 FreeSans 224 90 0 0 NN4BEG[8]
port 90 nsew signal tristate
flabel metal2 s 17682 9840 17738 10000 0 FreeSans 224 90 0 0 NN4BEG[9]
port 91 nsew signal tristate
flabel metal2 s 20258 9840 20314 10000 0 FreeSans 224 90 0 0 S1END[0]
port 92 nsew signal input
flabel metal2 s 20626 9840 20682 10000 0 FreeSans 224 90 0 0 S1END[1]
port 93 nsew signal input
flabel metal2 s 20994 9840 21050 10000 0 FreeSans 224 90 0 0 S1END[2]
port 94 nsew signal input
flabel metal2 s 21362 9840 21418 10000 0 FreeSans 224 90 0 0 S1END[3]
port 95 nsew signal input
flabel metal2 s 21730 9840 21786 10000 0 FreeSans 224 90 0 0 S2END[0]
port 96 nsew signal input
flabel metal2 s 22098 9840 22154 10000 0 FreeSans 224 90 0 0 S2END[1]
port 97 nsew signal input
flabel metal2 s 22466 9840 22522 10000 0 FreeSans 224 90 0 0 S2END[2]
port 98 nsew signal input
flabel metal2 s 22834 9840 22890 10000 0 FreeSans 224 90 0 0 S2END[3]
port 99 nsew signal input
flabel metal2 s 23202 9840 23258 10000 0 FreeSans 224 90 0 0 S2END[4]
port 100 nsew signal input
flabel metal2 s 23570 9840 23626 10000 0 FreeSans 224 90 0 0 S2END[5]
port 101 nsew signal input
flabel metal2 s 23938 9840 23994 10000 0 FreeSans 224 90 0 0 S2END[6]
port 102 nsew signal input
flabel metal2 s 24306 9840 24362 10000 0 FreeSans 224 90 0 0 S2END[7]
port 103 nsew signal input
flabel metal2 s 24674 9840 24730 10000 0 FreeSans 224 90 0 0 S2MID[0]
port 104 nsew signal input
flabel metal2 s 25042 9840 25098 10000 0 FreeSans 224 90 0 0 S2MID[1]
port 105 nsew signal input
flabel metal2 s 25410 9840 25466 10000 0 FreeSans 224 90 0 0 S2MID[2]
port 106 nsew signal input
flabel metal2 s 25778 9840 25834 10000 0 FreeSans 224 90 0 0 S2MID[3]
port 107 nsew signal input
flabel metal2 s 26146 9840 26202 10000 0 FreeSans 224 90 0 0 S2MID[4]
port 108 nsew signal input
flabel metal2 s 26514 9840 26570 10000 0 FreeSans 224 90 0 0 S2MID[5]
port 109 nsew signal input
flabel metal2 s 26882 9840 26938 10000 0 FreeSans 224 90 0 0 S2MID[6]
port 110 nsew signal input
flabel metal2 s 27250 9840 27306 10000 0 FreeSans 224 90 0 0 S2MID[7]
port 111 nsew signal input
flabel metal2 s 27618 9840 27674 10000 0 FreeSans 224 90 0 0 S4END[0]
port 112 nsew signal input
flabel metal2 s 31298 9840 31354 10000 0 FreeSans 224 90 0 0 S4END[10]
port 113 nsew signal input
flabel metal2 s 31666 9840 31722 10000 0 FreeSans 224 90 0 0 S4END[11]
port 114 nsew signal input
flabel metal2 s 32034 9840 32090 10000 0 FreeSans 224 90 0 0 S4END[12]
port 115 nsew signal input
flabel metal2 s 32402 9840 32458 10000 0 FreeSans 224 90 0 0 S4END[13]
port 116 nsew signal input
flabel metal2 s 32770 9840 32826 10000 0 FreeSans 224 90 0 0 S4END[14]
port 117 nsew signal input
flabel metal2 s 33138 9840 33194 10000 0 FreeSans 224 90 0 0 S4END[15]
port 118 nsew signal input
flabel metal2 s 27986 9840 28042 10000 0 FreeSans 224 90 0 0 S4END[1]
port 119 nsew signal input
flabel metal2 s 28354 9840 28410 10000 0 FreeSans 224 90 0 0 S4END[2]
port 120 nsew signal input
flabel metal2 s 28722 9840 28778 10000 0 FreeSans 224 90 0 0 S4END[3]
port 121 nsew signal input
flabel metal2 s 29090 9840 29146 10000 0 FreeSans 224 90 0 0 S4END[4]
port 122 nsew signal input
flabel metal2 s 29458 9840 29514 10000 0 FreeSans 224 90 0 0 S4END[5]
port 123 nsew signal input
flabel metal2 s 29826 9840 29882 10000 0 FreeSans 224 90 0 0 S4END[6]
port 124 nsew signal input
flabel metal2 s 30194 9840 30250 10000 0 FreeSans 224 90 0 0 S4END[7]
port 125 nsew signal input
flabel metal2 s 30562 9840 30618 10000 0 FreeSans 224 90 0 0 S4END[8]
port 126 nsew signal input
flabel metal2 s 30930 9840 30986 10000 0 FreeSans 224 90 0 0 S4END[9]
port 127 nsew signal input
flabel metal2 s 33506 9840 33562 10000 0 FreeSans 224 90 0 0 SS4END[0]
port 128 nsew signal input
flabel metal2 s 37186 9840 37242 10000 0 FreeSans 224 90 0 0 SS4END[10]
port 129 nsew signal input
flabel metal2 s 37554 9840 37610 10000 0 FreeSans 224 90 0 0 SS4END[11]
port 130 nsew signal input
flabel metal2 s 37922 9840 37978 10000 0 FreeSans 224 90 0 0 SS4END[12]
port 131 nsew signal input
flabel metal2 s 38290 9840 38346 10000 0 FreeSans 224 90 0 0 SS4END[13]
port 132 nsew signal input
flabel metal2 s 38658 9840 38714 10000 0 FreeSans 224 90 0 0 SS4END[14]
port 133 nsew signal input
flabel metal2 s 39026 9840 39082 10000 0 FreeSans 224 90 0 0 SS4END[15]
port 134 nsew signal input
flabel metal2 s 33874 9840 33930 10000 0 FreeSans 224 90 0 0 SS4END[1]
port 135 nsew signal input
flabel metal2 s 34242 9840 34298 10000 0 FreeSans 224 90 0 0 SS4END[2]
port 136 nsew signal input
flabel metal2 s 34610 9840 34666 10000 0 FreeSans 224 90 0 0 SS4END[3]
port 137 nsew signal input
flabel metal2 s 34978 9840 35034 10000 0 FreeSans 224 90 0 0 SS4END[4]
port 138 nsew signal input
flabel metal2 s 35346 9840 35402 10000 0 FreeSans 224 90 0 0 SS4END[5]
port 139 nsew signal input
flabel metal2 s 35714 9840 35770 10000 0 FreeSans 224 90 0 0 SS4END[6]
port 140 nsew signal input
flabel metal2 s 36082 9840 36138 10000 0 FreeSans 224 90 0 0 SS4END[7]
port 141 nsew signal input
flabel metal2 s 36450 9840 36506 10000 0 FreeSans 224 90 0 0 SS4END[8]
port 142 nsew signal input
flabel metal2 s 36818 9840 36874 10000 0 FreeSans 224 90 0 0 SS4END[9]
port 143 nsew signal input
flabel metal2 s 1858 0 1914 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 39394 9840 39450 10000 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6659 1040 6979 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 18089 1040 18409 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 29519 1040 29839 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 40949 1040 41269 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 12374 1040 12694 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 23804 1040 24124 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 35234 1040 35554 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 46664 1040 46984 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 23966 8160 23966 8160 0 vccd1
rlabel via1 24044 8704 24044 8704 0 vssd1
rlabel metal2 4147 68 4147 68 0 FrameStrobe[0]
rlabel metal2 26174 415 26174 415 0 FrameStrobe[10]
rlabel metal2 28435 68 28435 68 0 FrameStrobe[11]
rlabel metal2 30643 68 30643 68 0 FrameStrobe[12]
rlabel metal2 32851 68 32851 68 0 FrameStrobe[13]
rlabel metal2 35059 68 35059 68 0 FrameStrobe[14]
rlabel metal2 37267 68 37267 68 0 FrameStrobe[15]
rlabel metal2 39475 68 39475 68 0 FrameStrobe[16]
rlabel metal2 41683 68 41683 68 0 FrameStrobe[17]
rlabel metal2 43891 68 43891 68 0 FrameStrobe[18]
rlabel metal2 46191 68 46191 68 0 FrameStrobe[19]
rlabel metal2 6355 68 6355 68 0 FrameStrobe[1]
rlabel metal2 8563 68 8563 68 0 FrameStrobe[2]
rlabel metal2 10771 68 10771 68 0 FrameStrobe[3]
rlabel metal2 12979 68 12979 68 0 FrameStrobe[4]
rlabel metal2 15187 68 15187 68 0 FrameStrobe[5]
rlabel metal2 17395 68 17395 68 0 FrameStrobe[6]
rlabel metal2 19603 68 19603 68 0 FrameStrobe[7]
rlabel metal2 21811 68 21811 68 0 FrameStrobe[8]
rlabel metal2 24111 68 24111 68 0 FrameStrobe[9]
rlabel metal2 39790 9190 39790 9190 0 FrameStrobe_O[0]
rlabel metal2 43470 9836 43470 9836 0 FrameStrobe_O[10]
rlabel metal2 43838 9836 43838 9836 0 FrameStrobe_O[11]
rlabel metal2 44206 9836 44206 9836 0 FrameStrobe_O[12]
rlabel metal2 44574 8680 44574 8680 0 FrameStrobe_O[13]
rlabel metal2 44942 8340 44942 8340 0 FrameStrobe_O[14]
rlabel metal1 45080 7446 45080 7446 0 FrameStrobe_O[15]
rlabel metal2 45678 8680 45678 8680 0 FrameStrobe_O[16]
rlabel metal1 46138 6970 46138 6970 0 FrameStrobe_O[17]
rlabel metal2 46414 8680 46414 8680 0 FrameStrobe_O[18]
rlabel metal1 46276 8058 46276 8058 0 FrameStrobe_O[19]
rlabel metal1 40664 8330 40664 8330 0 FrameStrobe_O[1]
rlabel metal1 40848 8058 40848 8058 0 FrameStrobe_O[2]
rlabel metal2 40894 9224 40894 9224 0 FrameStrobe_O[3]
rlabel metal2 41262 9190 41262 9190 0 FrameStrobe_O[4]
rlabel metal2 41630 9088 41630 9088 0 FrameStrobe_O[5]
rlabel metal2 41998 9122 41998 9122 0 FrameStrobe_O[6]
rlabel metal2 42366 9836 42366 9836 0 FrameStrobe_O[7]
rlabel metal2 42734 9224 42734 9224 0 FrameStrobe_O[8]
rlabel metal2 43102 9836 43102 9836 0 FrameStrobe_O[9]
rlabel metal1 23920 1734 23920 1734 0 FrameStrobe_O_i\[0\]
rlabel metal1 27370 2074 27370 2074 0 FrameStrobe_O_i\[10\]
rlabel metal1 29532 2074 29532 2074 0 FrameStrobe_O_i\[11\]
rlabel metal2 31418 2244 31418 2244 0 FrameStrobe_O_i\[12\]
rlabel metal1 33948 2074 33948 2074 0 FrameStrobe_O_i\[13\]
rlabel metal1 36110 2074 36110 2074 0 FrameStrobe_O_i\[14\]
rlabel metal1 38318 2074 38318 2074 0 FrameStrobe_O_i\[15\]
rlabel metal1 44666 2074 44666 2074 0 FrameStrobe_O_i\[16\]
rlabel metal1 42872 2074 42872 2074 0 FrameStrobe_O_i\[17\]
rlabel metal2 44758 2074 44758 2074 0 FrameStrobe_O_i\[18\]
rlabel metal1 45908 2074 45908 2074 0 FrameStrobe_O_i\[19\]
rlabel metal1 23460 1802 23460 1802 0 FrameStrobe_O_i\[1\]
rlabel metal1 23460 2074 23460 2074 0 FrameStrobe_O_i\[2\]
rlabel metal1 24288 2074 24288 2074 0 FrameStrobe_O_i\[3\]
rlabel metal1 23644 1530 23644 1530 0 FrameStrobe_O_i\[4\]
rlabel metal1 23736 1462 23736 1462 0 FrameStrobe_O_i\[5\]
rlabel metal2 22402 2244 22402 2244 0 FrameStrobe_O_i\[6\]
rlabel metal1 20700 2074 20700 2074 0 FrameStrobe_O_i\[7\]
rlabel metal1 22954 2074 22954 2074 0 FrameStrobe_O_i\[8\]
rlabel metal1 25070 2074 25070 2074 0 FrameStrobe_O_i\[9\]
rlabel metal2 1150 8952 1150 8952 0 N1BEG[0]
rlabel metal2 1518 8680 1518 8680 0 N1BEG[1]
rlabel metal1 2438 7956 2438 7956 0 N1BEG[2]
rlabel metal1 2024 8602 2024 8602 0 N1BEG[3]
rlabel metal1 2162 8364 2162 8364 0 N2BEG[0]
rlabel metal2 2990 9224 2990 9224 0 N2BEG[1]
rlabel metal1 3220 8602 3220 8602 0 N2BEG[2]
rlabel metal1 3588 8602 3588 8602 0 N2BEG[3]
rlabel metal2 4094 8952 4094 8952 0 N2BEG[4]
rlabel metal1 4232 8602 4232 8602 0 N2BEG[5]
rlabel metal1 4738 8058 4738 8058 0 N2BEG[6]
rlabel metal1 4738 8602 4738 8602 0 N2BEG[7]
rlabel metal1 5290 8602 5290 8602 0 N2BEGb[0]
rlabel metal1 5796 8602 5796 8602 0 N2BEGb[1]
rlabel metal1 6164 8602 6164 8602 0 N2BEGb[2]
rlabel metal2 6670 9309 6670 9309 0 N2BEGb[3]
rlabel metal2 6762 9231 6762 9231 0 N2BEGb[4]
rlabel metal1 7314 8058 7314 8058 0 N2BEGb[5]
rlabel metal1 7452 8602 7452 8602 0 N2BEGb[6]
rlabel metal1 7682 8330 7682 8330 0 N2BEGb[7]
rlabel metal1 8142 8602 8142 8602 0 N4BEG[0]
rlabel metal1 11960 8602 11960 8602 0 N4BEG[10]
rlabel metal2 12558 9785 12558 9785 0 N4BEG[11]
rlabel metal1 12788 8058 12788 8058 0 N4BEG[12]
rlabel metal1 13064 8602 13064 8602 0 N4BEG[13]
rlabel metal1 13340 8330 13340 8330 0 N4BEG[14]
rlabel metal1 13892 8602 13892 8602 0 N4BEG[15]
rlabel metal1 8970 8602 8970 8602 0 N4BEG[1]
rlabel metal2 9246 8952 9246 8952 0 N4BEG[2]
rlabel metal1 8602 8568 8602 8568 0 N4BEG[3]
rlabel metal1 9522 8534 9522 8534 0 N4BEG[4]
rlabel metal1 10212 8058 10212 8058 0 N4BEG[5]
rlabel metal1 10258 8602 10258 8602 0 N4BEG[6]
rlabel metal1 10810 8602 10810 8602 0 N4BEG[7]
rlabel metal1 11316 8602 11316 8602 0 N4BEG[8]
rlabel metal2 11822 8952 11822 8952 0 N4BEG[9]
rlabel metal2 14398 8952 14398 8952 0 NN4BEG[0]
rlabel metal2 18078 9224 18078 9224 0 NN4BEG[10]
rlabel metal1 18538 8602 18538 8602 0 NN4BEG[11]
rlabel metal1 18906 8602 18906 8602 0 NN4BEG[12]
rlabel metal2 19182 9445 19182 9445 0 NN4BEG[13]
rlabel metal1 20562 8364 20562 8364 0 NN4BEG[14]
rlabel metal1 20056 8602 20056 8602 0 NN4BEG[15]
rlabel metal1 14858 8058 14858 8058 0 NN4BEG[1]
rlabel metal1 14812 8602 14812 8602 0 NN4BEG[2]
rlabel metal1 15272 8602 15272 8602 0 NN4BEG[3]
rlabel metal1 15732 8058 15732 8058 0 NN4BEG[4]
rlabel metal1 16008 8602 16008 8602 0 NN4BEG[5]
rlabel metal1 16422 8602 16422 8602 0 NN4BEG[6]
rlabel metal1 17020 8058 17020 8058 0 NN4BEG[7]
rlabel metal1 17204 8602 17204 8602 0 NN4BEG[8]
rlabel metal1 17664 8602 17664 8602 0 NN4BEG[9]
rlabel metal2 20286 8612 20286 8612 0 S1END[0]
rlabel metal2 20654 9377 20654 9377 0 S1END[1]
rlabel metal2 21022 9241 21022 9241 0 S1END[2]
rlabel metal2 21390 9785 21390 9785 0 S1END[3]
rlabel metal2 21758 9190 21758 9190 0 S2END[0]
rlabel metal1 21758 8466 21758 8466 0 S2END[1]
rlabel metal2 22494 9700 22494 9700 0 S2END[2]
rlabel metal2 22862 9836 22862 9836 0 S2END[3]
rlabel metal2 23230 9836 23230 9836 0 S2END[4]
rlabel metal2 23598 9836 23598 9836 0 S2END[5]
rlabel metal2 23966 9836 23966 9836 0 S2END[6]
rlabel metal2 24334 9190 24334 9190 0 S2END[7]
rlabel metal2 24702 9836 24702 9836 0 S2MID[0]
rlabel metal2 25070 9836 25070 9836 0 S2MID[1]
rlabel metal2 25438 9836 25438 9836 0 S2MID[2]
rlabel metal2 25806 9836 25806 9836 0 S2MID[3]
rlabel metal2 26174 9836 26174 9836 0 S2MID[4]
rlabel metal2 26542 9836 26542 9836 0 S2MID[5]
rlabel metal2 26910 9836 26910 9836 0 S2MID[6]
rlabel metal2 27278 9836 27278 9836 0 S2MID[7]
rlabel metal2 27646 9836 27646 9836 0 S4END[0]
rlabel metal2 31326 9836 31326 9836 0 S4END[10]
rlabel metal2 31694 9156 31694 9156 0 S4END[11]
rlabel metal2 32062 9836 32062 9836 0 S4END[12]
rlabel metal2 32430 9836 32430 9836 0 S4END[13]
rlabel metal2 32798 9836 32798 9836 0 S4END[14]
rlabel metal2 33166 9836 33166 9836 0 S4END[15]
rlabel metal2 28014 9836 28014 9836 0 S4END[1]
rlabel metal2 28382 9836 28382 9836 0 S4END[2]
rlabel metal2 28750 9156 28750 9156 0 S4END[3]
rlabel metal2 29118 9836 29118 9836 0 S4END[4]
rlabel metal2 29486 9836 29486 9836 0 S4END[5]
rlabel metal2 29854 9836 29854 9836 0 S4END[6]
rlabel metal2 30222 9156 30222 9156 0 S4END[7]
rlabel metal2 30590 9224 30590 9224 0 S4END[8]
rlabel metal2 30958 9836 30958 9836 0 S4END[9]
rlabel metal2 33534 9836 33534 9836 0 SS4END[0]
rlabel metal2 37214 9156 37214 9156 0 SS4END[10]
rlabel metal2 37582 9836 37582 9836 0 SS4END[11]
rlabel metal2 37950 9836 37950 9836 0 SS4END[12]
rlabel metal2 38318 9836 38318 9836 0 SS4END[13]
rlabel metal2 38686 9836 38686 9836 0 SS4END[14]
rlabel metal2 39054 9836 39054 9836 0 SS4END[15]
rlabel metal2 33902 9836 33902 9836 0 SS4END[1]
rlabel metal2 34270 9156 34270 9156 0 SS4END[2]
rlabel metal2 34638 9836 34638 9836 0 SS4END[3]
rlabel metal2 35006 9156 35006 9156 0 SS4END[4]
rlabel metal2 35374 9836 35374 9836 0 SS4END[5]
rlabel metal2 35742 9156 35742 9156 0 SS4END[6]
rlabel metal2 36110 9836 36110 9836 0 SS4END[7]
rlabel metal2 36478 9836 36478 9836 0 SS4END[8]
rlabel metal2 36846 9836 36846 9836 0 SS4END[9]
rlabel metal2 1939 68 1939 68 0 UserCLK
rlabel metal2 39422 9224 39422 9224 0 UserCLKo
rlabel metal1 4370 1224 4370 1224 0 net1
rlabel metal1 44344 1530 44344 1530 0 net10
rlabel metal2 3266 7667 3266 7667 0 net100
rlabel metal2 6486 7344 6486 7344 0 net101
rlabel metal2 4370 7106 4370 7106 0 net102
rlabel metal2 8326 7259 8326 7259 0 net103
rlabel metal2 20746 6868 20746 6868 0 net104
rlabel metal2 9706 7718 9706 7718 0 net105
rlabel metal2 12742 9622 12742 9622 0 net106
rlabel metal2 13662 9146 13662 9146 0 net107
rlabel metal1 17158 9826 17158 9826 0 net108
rlabel metal2 16514 7004 16514 7004 0 net109
rlabel metal1 45908 1530 45908 1530 0 net11
rlabel metal1 21620 8058 21620 8058 0 net110
rlabel metal2 18170 7735 18170 7735 0 net111
rlabel metal2 21298 8755 21298 8755 0 net112
rlabel metal1 20976 8058 20976 8058 0 net113
rlabel metal1 8142 8432 8142 8432 0 net114
rlabel metal1 28244 7718 28244 7718 0 net115
rlabel metal1 28658 8058 28658 8058 0 net116
rlabel metal2 13754 8381 13754 8381 0 net117
rlabel metal2 20930 9741 20930 9741 0 net118
rlabel metal1 13386 8908 13386 8908 0 net119
rlabel metal1 6578 816 6578 816 0 net12
rlabel metal2 27094 8874 27094 8874 0 net120
rlabel metal1 23644 8058 23644 8058 0 net121
rlabel metal1 17066 9928 17066 9928 0 net122
rlabel metal2 21390 8993 21390 8993 0 net123
rlabel metal2 21666 9435 21666 9435 0 net124
rlabel metal1 15962 8024 15962 8024 0 net125
rlabel via2 21666 9027 21666 9027 0 net126
rlabel via2 14858 8517 14858 8517 0 net127
rlabel metal1 13570 8432 13570 8432 0 net128
rlabel metal1 14582 7820 14582 7820 0 net129
rlabel metal2 19918 1428 19918 1428 0 net13
rlabel metal1 20930 7412 20930 7412 0 net130
rlabel metal1 18032 8058 18032 8058 0 net131
rlabel metal1 18400 8058 18400 8058 0 net132
rlabel metal2 18814 8262 18814 8262 0 net133
rlabel metal1 19642 7242 19642 7242 0 net134
rlabel metal2 20194 7990 20194 7990 0 net135
rlabel metal1 19964 8058 19964 8058 0 net136
rlabel metal1 20562 7888 20562 7888 0 net137
rlabel metal1 19734 7344 19734 7344 0 net138
rlabel metal2 22954 7276 22954 7276 0 net139
rlabel metal2 23322 1292 23322 1292 0 net14
rlabel metal1 15778 6936 15778 6936 0 net140
rlabel metal2 21482 8908 21482 8908 0 net141
rlabel metal2 21206 7140 21206 7140 0 net142
rlabel metal2 17250 8092 17250 8092 0 net143
rlabel metal1 20654 8058 20654 8058 0 net144
rlabel metal1 17756 8058 17756 8058 0 net145
rlabel metal1 25346 1734 25346 1734 0 net146
rlabel metal1 21206 952 21206 952 0 net15
rlabel metal1 23230 918 23230 918 0 net16
rlabel metal1 19274 1190 19274 1190 0 net17
rlabel metal1 19964 1530 19964 1530 0 net18
rlabel metal1 22264 1530 22264 1530 0 net19
rlabel metal1 26726 1530 26726 1530 0 net2
rlabel metal1 24380 1530 24380 1530 0 net20
rlabel metal1 20056 7174 20056 7174 0 net21
rlabel metal2 19550 7956 19550 7956 0 net22
rlabel metal1 20516 7514 20516 7514 0 net23
rlabel metal1 20700 7854 20700 7854 0 net24
rlabel metal2 21206 8058 21206 8058 0 net25
rlabel metal2 21482 8058 21482 8058 0 net26
rlabel metal1 21804 7854 21804 7854 0 net27
rlabel metal2 22034 8058 22034 8058 0 net28
rlabel metal1 22678 7378 22678 7378 0 net29
rlabel metal1 28888 1530 28888 1530 0 net3
rlabel metal1 22310 7820 22310 7820 0 net30
rlabel metal1 22586 7888 22586 7888 0 net31
rlabel metal1 23506 7854 23506 7854 0 net32
rlabel metal1 24242 7412 24242 7412 0 net33
rlabel metal1 24242 7888 24242 7888 0 net34
rlabel metal1 25116 7854 25116 7854 0 net35
rlabel metal1 25346 7888 25346 7888 0 net36
rlabel metal2 26174 8092 26174 8092 0 net37
rlabel metal1 26542 7854 26542 7854 0 net38
rlabel metal1 26772 7854 26772 7854 0 net39
rlabel metal1 31050 1530 31050 1530 0 net4
rlabel metal1 27094 7854 27094 7854 0 net40
rlabel metal1 27370 7854 27370 7854 0 net41
rlabel metal1 28152 7378 28152 7378 0 net42
rlabel metal1 24886 7480 24886 7480 0 net43
rlabel metal2 32154 8840 32154 8840 0 net44
rlabel metal1 32522 8500 32522 8500 0 net45
rlabel metal2 29026 7922 29026 7922 0 net46
rlabel metal2 33258 9078 33258 9078 0 net47
rlabel metal2 27554 8058 27554 8058 0 net48
rlabel metal1 28060 7854 28060 7854 0 net49
rlabel metal1 33304 1530 33304 1530 0 net5
rlabel metal1 28428 7854 28428 7854 0 net50
rlabel metal1 28658 7888 28658 7888 0 net51
rlabel metal1 29164 7854 29164 7854 0 net52
rlabel metal1 29394 7888 29394 7888 0 net53
rlabel metal1 30084 7854 30084 7854 0 net54
rlabel metal1 25714 7854 25714 7854 0 net55
rlabel metal1 25944 7854 25944 7854 0 net56
rlabel metal2 33626 9044 33626 9044 0 net57
rlabel metal1 37168 8262 37168 8262 0 net58
rlabel metal2 37674 8942 37674 8942 0 net59
rlabel metal1 35420 1530 35420 1530 0 net6
rlabel metal2 36938 7922 36938 7922 0 net60
rlabel metal2 37122 8058 37122 8058 0 net61
rlabel metal2 38778 7871 38778 7871 0 net62
rlabel metal2 39146 8908 39146 8908 0 net63
rlabel metal2 33994 8874 33994 8874 0 net64
rlabel metal1 33672 8330 33672 8330 0 net65
rlabel metal1 34408 8602 34408 8602 0 net66
rlabel metal2 35098 8211 35098 8211 0 net67
rlabel metal1 35282 8602 35282 8602 0 net68
rlabel metal2 35834 8143 35834 8143 0 net69
rlabel metal1 37628 1530 37628 1530 0 net7
rlabel metal2 36202 8738 36202 8738 0 net70
rlabel metal2 36570 8806 36570 8806 0 net71
rlabel metal1 36708 8330 36708 8330 0 net72
rlabel metal2 2162 1088 2162 1088 0 net73
rlabel metal1 25254 2516 25254 2516 0 net74
rlabel metal2 45126 6290 45126 6290 0 net75
rlabel metal2 44022 5644 44022 5644 0 net76
rlabel metal1 41078 9078 41078 9078 0 net77
rlabel metal1 40756 7310 40756 7310 0 net78
rlabel metal1 42826 2584 42826 2584 0 net79
rlabel metal2 44114 1564 44114 1564 0 net8
rlabel metal1 43056 7378 43056 7378 0 net80
rlabel metal1 45402 2618 45402 2618 0 net81
rlabel metal1 43838 2618 43838 2618 0 net82
rlabel metal1 45908 7378 45908 7378 0 net83
rlabel metal2 45770 4759 45770 4759 0 net84
rlabel metal1 24886 2312 24886 2312 0 net85
rlabel metal1 40526 7854 40526 7854 0 net86
rlabel metal1 41262 8466 41262 8466 0 net87
rlabel metal1 41538 8432 41538 8432 0 net88
rlabel metal1 24472 1734 24472 1734 0 net89
rlabel metal1 42182 1530 42182 1530 0 net9
rlabel metal2 36110 5235 36110 5235 0 net90
rlabel metal1 21206 2040 21206 2040 0 net91
rlabel metal2 24978 2397 24978 2397 0 net92
rlabel metal1 40986 9010 40986 9010 0 net93
rlabel metal1 2162 7480 2162 7480 0 net94
rlabel metal2 20010 7616 20010 7616 0 net95
rlabel metal1 2622 7786 2622 7786 0 net96
rlabel metal1 1978 8976 1978 8976 0 net97
rlabel metal2 2346 8143 2346 8143 0 net98
rlabel metal1 13570 9316 13570 9316 0 net99
<< properties >>
string FIXED_BBOX 0 0 48000 10000
<< end >>
